ELF              ؗ4   �     4    (      4   4�4��   �            �   ��                    � �H� H�          `� `�`�0  �b          0 0�0��   �              ��              /lib/ld-linux.so.2           GNU              a   g   R      C   6       	       +   I   5          G   ?           ^   c   4      J   A      0              M   Z       X   B   [   V   _       U   2   Y           #       a          W   7   K   d              /   F       e   <   %           S       9           `       T             )      .   O                      (       *   b                   f      !       ]       H                                                                                                                                                                                      &                   $      ,       '         3       -          ;   
      "                           8              D   >         N              L      P           =       @   1                 \   Q       E       :                   	  H�:         X�&      E   h��     �   x�Y,     )  ��?     �   ���      �  ��g     �   ��1     J  Ȓm        ؒ      M   0�     ���  �q      V   ���     �  �|        �8      �  (�2      5  8�%      V  H�q      /  X�:     �  h�#        x�Z        ��     �  ��6      �  ���      j  ���      �  ȓ6      �  ؓL      \  �_     <  ��$     6  �x      �  �9      �  (��      /  8�|     C  H�{      �  X�:      ^    �     
 O  h��       x�#      w  ��6      d   ��<      V  ��e      �  ��:      q   Ȕ[      �   ��     f  ��     �  ؔ&     �  �     �  ��'      #  �@      #  �S       (�F     d  8�       H�U     �  X��      m  h��      �   x�2      |  ���        ��     ���  ���      �  ���     �  ���        ȕ+      �   ؕ0      <  �C      ~   h2      q  ��|      U  ��     �   �      I  (��      �   8�|      �  H��      �  X��       h�4        ��     ���   �     ��  x��      '  ��     ��]  ��5         ���      (  ��C      �  ��      �  ��     �  Ȗ�      �  ؖ5      E  �6      �  �2       ���      �  �:      �   �4      �  (�q     �  8�N      �   H�u         X�&        h��                     s  x�q      �  ��|      �   ���      �   ��C      �  ���      ,               �   ȗ0       libm.so.6 sin tan acos _Jv_RegisterClasses __gmon_start__ libz.so.1 deflate _DYNAMIC inflate _init inflateInit_ deflateInit_ _fini _GLOBAL_OFFSET_TABLE_ inflateEnd deflateEnd libc.so.6 strcpy asctime __strtod_internal stdout vsprintf fdopen geteuid xdrmem_create getenv getpid qsort fscanf fgets execl perror creat getuid system feof malloc remove isatty sleep fflush lseek pipe xdr_double __ctype_tolower_loc calloc fprintf kill strcat dcgettext fseek stdin wait umask signal read strncmp strncpy unlink realloc _IO_getc strtok fork sscanf localtime memset ftell strcmp getpwuid dup gethostname fclose setlocale stderr fputc __ctype_b_loc fwrite access __xstat rewind xdr_float __errno_location bindtextdomain fopen fileno _IO_stdin_used _exit __libc_start_main strchr fputs mkdir free _edata __bss_start _end GLIBC_2.0 GLIBC_2.3 GLIBC_2.1                                                                                                                             ii   ,        �          ii   6     ii   @     ii   ,      ��e  ��,  ��-  ��R  (�  ,�  0�  4�  8�  <�  @�  D�  H�	  L�
  P�  T�  X�  \�  `�  d�  h�  l�  p�  t�  x�  |�  ��  ��  ��  ��  ��  ��  ��  ��  ��   ��!  ��"  ��#  ��%  ��&  ��'  ��(  ��)  Ē*  Ȓ+  ̒.  В/  Ԓ0  ؒ1  ܒ2  ��3  �4  �5  �6  �7  ��8  ��9  ��;   �<  �=  �>  �?  �@  �B  �C  �D   �E  $�F  (�G  ,�H  0�I  4�L  8�N  <�O  @�P  D�Q  H�S  L�T  P�U  T�W  X�X  \�Y  `�Z  d�[  h�\  l�]  p�^  t�`  x�a  |�b  ��c  ��d  ��f  U�����  �,  �� �� �5 ��%$�    �%(�h    ������%,�h   ������%0�h   ������%4�h   �����%8�h    �����%<�h(   �����%@�h0   �����%D�h8   �p����%H�h@   �`����%L�hH   �P����%P�hP   �@����%T�hX   �0����%X�h`   � ����%\�hh   �����%`�hp   � ����%d�hx   ������%h�h�   ������%l�h�   ������%p�h�   ������%t�h�   �����%x�h�   �����%|�h�   �����%��h�   �����%��h�   �p����%��h�   �`����%��h�   �P����%��h�   �@����%��h�   �0����%��h�   � ����%��h�   �����%��h�   � ����%��h�   ������%��h   ������%��h  ������%��h  ������%��h  �����%��h   �����%��h(  �����%��h0  �����%Ēh8  �p����%Ȓh@  �`����%̒hH  �P����%ВhP  �@����%ԒhX  �0����%ؒh`  � ����%ܒhh  �����%��hp  � ����%�hx  ������%�h�  ������%�h�  ������%�h�  ������%��h�  �����%��h�  �����%��h�  �����% �h�  �����%�h�  �p����%�h�  �`����%�h�  �P����%�h�  �@����%�h�  �0����%�h�  � ����%�h�  �����% �h�  � ����%$�h�  ������%(�h   ������%,�h  ������%0�h  ������%4�h  �����%8�h   �����%<�h(  �����%@�h0  �����%D�h8  �p����%H�h@  �`����%L�hH  �P����%P�hP  �@����%T�hX  �0����%X�h`  � ����%\�hh  �����%`�hp  � ����%d�hx  ������%h�h�  ������%l�h�  ������%p�h�  ������%t�h�  �����%x�h�  �����%|�h�  �����%��h�  �����%��h�  �p����%��h�  �`���1�^����PTRh2h�1QVh���������U��SP�    [��� ��p  ��t�Ћ]��Ð�U����=�� u)�h����t�����h��ҡh����u�����É�U�������t�    ��t��h��g�����Ð�U��WVS��|  ������]�3ǅ����    �.  �m_  � �2�~^  � �5�@   �@    �@�5�@,�5�������Q^  � `6�@   �@   �@�5�������+^  � �5�@   �@    �@s6�� ����^  � �5�@   �@    �@�5�������]  �  6�@   �@    �@6������]  � 6�@   �@    �@ 3������]  �  W�@   �@!6�@    �@    �@`3������\  � q�@#6���\  � p�@)6��XZS�u�7^  ����t��j�  ����j ��  �$C6�Z��������1��~ ��������������Ph�s������p�	�����������Ph�O�������p�������Ht��hQ6�  ��� ����B���  P������Ph�O�r������Ht��hd6�c  �(7܍����݅����������Eu��h�3�;  ������B����  P������Ph�O�rǅ����    �G�����Ht��h�6��  ������B���R  V������Ph�O�r������Ht��h�3�  �v ������@�w��������������t
ǅ����   ����������  �������p����  Sh�6Vh�6�  ��������  ��h ��)  XZS�������p���  �������J  ��������Ph �������������j R���  �������������� ��u��h 4��  ��������tW������h�6�5�����������������������
  �����������$�6  ��������  ǅ����    ������9�����}H݅����1ҋ�����@P���$���������\�D    �D    �    ��9ȉ�����|����  H~��h`4�  ����������t�5��j$jh�4���������������ǅ����    �  ǅ����    ǅ����    ������9�������  1�������9������z  �������������0�D0���,���l����������ݝ�����0����D0�l��݅���������󋍘������07�R  �����������������������������$ݝx����	  �� ��݅x����  ��ܵ����ٽ����f������%����   f������٭������٭����ٽ����ݝ����f�������f������݅����٭����۝����٭�����������X�;�������  ����    �D݅���������������U  ��������������  ���؋������D0�������l���D��\�v ��������������9������Y�����������tPj��������������y  ��������������������9������������������~.��1ҋ������D������E�  ������\��Ku��؋�������tPjjj�y  ������������������������tj��������t�5��j$jh�4�C�����������������������W�  ����������tQjjj�y  ����W�S����$    ������������~�1��������D7����������Eu'P�47�t7�t7�t7�t7h�6�5��������� ��Ku���������ɍ����Q�B����������um����������u$�������D0�������l���B�A�Z�*�����������������h�6�����S� ����$�  ǅ����   �����������������k����؃�h�6��G  ����������������h 5��PVh�6�����S�����$��QVh7���������Ph �R������j �5��������h`5�ǅ����    ǅ����    �����ǅ����   �����(7܍����ݝ����������U��WVS�������1��ы}����ЍP�1�9��E�    �E�    }'��u�}�<7/�  �E܋E�9��؉��E�9U�|ھ����1҈Ћ}�����щM؋}�����ҋu؍D�ËE����P�Y  �E�    �}��9}�E�},C�v ��S�7  �U�M���������  �E�u�9u�|؋}�O�E�    9}��E�    �}���   �]��v ���u�3������1������������֋E�~������}�u �}�E��M���M܈G�u܋u��}��}�M�9</t(��t$�u܈�E�F�u܋}�U�:</t��t��ދ�M܃�� �u�3�P����E�u��E����9u��P������}��u�E��4��4����M��������1��ى������H�E܋]�u���</t9��t5�]܈�E�C�]܋u�}�7��/��tF��t�}�M����ԋE�M����}�� ���u�E�U��4������E�M��E��e�[^_�Ë]�u������E��E�    ������5��jjh`7������$������������U��WVS��  �E1�����  ��P������S��  �$��  �������� ��  Sh�7h�7������V�\�����h�7h�7������P�C���XZhzz�5H�������������c  ��h�qV������������H  �������v PSh   V���������tV������<cu	������dt�<pu������lu	������ot��t���WV�������밃�������PPP�uW������� 떃�S�}����<$�u���Y�5H��)���XZhzz�5���'���������t~��h�q������P�
���������ta�PSh   V�3�������t��WV�2������݃�S�����<$�����Y�5������Z�5������X�5H������e�[^_�Ã�h�7�g
  �$�����<$��������h�7�H
  �$�����<$�����QSh�7������V������S�2�����U��E���   �EP�]���  �E��E����m����m��������������]��E��u��}�f�E�%����   f�E��m����m��}��]�f�E��f�E��E��m��]��m��E�@�Ð��U���E�E����� 8����������E���E���8  �����������Eu����v �������������	  �������������t�����������E����   ������������Eu����v ��������������   �������������t�����������E����   ������������Eu����v ����������ua�v ������������t�����������Eu������������Eu/����������������u������u	�   �É�1����������������������\������2������������������U��WVS��  ���  ��h�qP����4����������  PjjhC9�h����E����~$1��]��E�D0����������E��  ��Ku��W������  [^h�qP�H��������������  h�xhO9��d���P�5�������Ƌ�d���1�H��9��  WjjhT9�����Wj!jh 8������ Wj
jhd9����Wjjho9������ �}d��9��9P��d����t��h`8W����XZhtdj"j"h�=h�8��h���V�B�����W�)���_X��h���P������S������5H��5��h�9S������S�t�  �]����t*�M��t9Rjjj�o  �5��j$jh�8������� �E��t���uV�	������e�[^1�_��Q�4�h�OW�������d���CH��9�|�������P�E�40�t0�t0�t0�t0h�6W������ �2�����h 9�  �U����E��~��P��������t
�Ð�   ���h�9�  U����U�ҋE~ ��~��PR�B�������t�Ð�   �吺   �ك�h�9�<  U����U�ҋE~$��t��RP�N�������t�Ð��R������됺   �Ճ�h�9��  U�����������U������    ���  �?��o  �����t7��q  �����������u1����    ���  �?�Ð�   ������E�P�E�P�0  �u��u��u��u��  �   ��U����=���E�E�E�E t%���������������������]��E�����Ív �� �\$�\$�\$�$�y  ��v U��VS��`�E�]ЍE��EP�]ȍE��EP�]��E��E(P�]��E��E0P�]��E8���]��E@�$�u��u��u��u��]��] �u$�u��u�VS�u��u��u��u��u��u��  ��P����~
�e�[^�Ív ��VS�u��u��u��u��u��u��u��u��u��u��   �� �\$VS�u��u��u��u��u��u��u��u��u��u��m   ��0�$�u��u��u��u��u��u��u��u�VS�u��u��B   �� �\$�u��u��u��u��u��u��u��u��u��u��u��u��   ��0�$�[  �8�����U��S��t�E�E���]��]��E�E ���]��]��E0�E(���]��E������]��E��e��]�����������E��@�]���  �E�������E��@��  ���u��u���  XZ�u��u��]��  �E���������E�T  �E��E��E��E����u��������EȍE�P�E�P�E�P�E�P�u��u��u��u��u��u��u��u����\$�$�u��u��u��u���  ��P������   �E�������������u��������tT�u��u��u��u��u��u��u��u��������\$�u��u��u��u��u��u��u��u�������� �$�,  �]��Ív �u��u��u��u��u��u��u��u�������ِ����5��j3jh :�������u��u��u��u��u��u��u��u��u��u��u��u�Sh`:�5���������:��E��E��E��E����u��������E��������v �u��u��u��u��u��u��u��u��_����v ���0����U���E��������Eu���Ív U��VS���E�]�u�]��u$�u �u�u�#   ���]VS�u��u��   �]���e�[^����U���E�E������Eu���É�����U��S��  �EP�u������S����XZjS�   �$   �����U��S��  �����t1��]��ÐR�EP�u������S����YXj S�Z   ��U��U�������ÐU��1��=�� ��1҃} �����U��E���1��ÐU�����    1��Ív U��WVS�������tq�����uX�U��QtHPh�:h�:�@  ��Ph�:�5����������uh�O�5�������������e�[^_�ÐPh�:붃��u�u���ݍv ���u�u���   �H  ��������+  P�E���  Ph�:h�:�  ��Ph�:�5���L����}������   ��h�:h�:�x  ���1���������ӋE���]��E�u��}��SVW�5���  ����u���5�������$���������tI���5��j�����^�5���
����������t���    1��������j�b���������h�:��������ũ��u�u�  �׃�h�:�&���Ph�:��������u�u���U��WVS��(  j �����Y[h�O������W�����������XZhzzhn?�gf  ������t=VPh   W��������t����������t��<
��   B���u��S� g  ���  ����t��W������P�u�u�T   �� �<  ����t��t��SP�T�������u�e�[^1�_�Ív ��W������V�u�u�   �� �ؐ� �x���U��S���  �E��t�8 u�   �Ћ]��É�RPh�:�����S�����YXj S����������   u΃�hvS�a��������ú   t�Pj&jh�:�����f  PRh;h�:�
  ��Ph;S������ �{�  PPh;h�:��  ��Ph;S�����uPh;h�:��  ��Ph;S�e������EP�	�����PPh!;h�:�  ��Ph;S�6����E���ut@Ph';h�:�h  ��Ph;S������ Sj&jh�:�����$����1�����Ph.;�U��S��D��  ��t�8 u�   �]��Ð����  ��Ph7;�]�S�Z���XZh�qS��c  ������t4�E���ut.Ph�:h�:��  ��PhA;S�k����$�d  ��1��Qh�:��U��WVS���E� �U�E���1�< ��   <	��   <
��   1�����t < t<	t<
tB�G��t< t<	t<
u����   �E��D���E�u��K~9N��~���uj
N����������h�6�uhM;�u�����UB�U������uj ��������O��~���u�P������C��O���E��U��E��   �e�[^_�Ã��uj
�N���1����C<
t�< t�<	t�<
t�����F��U��WVS���  �]�; u1ҍe�[^��_��Q������P������VSƅ���� �8  ������   ����������W�X  ��1�@t���t�> uE1ې��S��  ������t���j RVW�u������P�3�  ��P�~����������k���C뾃�V��  ��1�@�S����> t���j PVW�u������P���  ��P�4��������!�����V��  ��������ߋu�A�����U��WVS��  �u�uV�u�����������tW������P������WV�+  ����u�e��[^_�É���WV�&�������U����������U������E�U�e�ȓ�̓����������������;���1��ÐU�����;�M�5�;�$���������������1���U���X��;�M�5�;�$���������������������������(7�������$�]��]�������E��$�]������YX�u��u��]�����XZ�u��u��]������E������E������E����Г���E����������������������������ؓ�����1��ÐU���X�E�e��;�5�;�(7�$�6�������������E����@u%������������ɀ�E��@�U���  ���������������������E��@u��������;�ȓ�]��E����������]�������������������E����@��t�E������ʀ�E��@�U��   �����������ɀ�E��@�U���   ���Г�E������ؓ����;�����M�����������;�����ȓ�E��E��������]�������;������������������������(7�m����������������������������������������m���������M��]�������؃��u��u��]��]�������E������]������E��������������������������v U��VS���E�]��E�]�] �u$�u�u�����XZVS�����E��]�E��]���e�[^������U��WVS��  �5��hR=h�6������S��  XZj S���������t+�E�    @�@�TXA�E� ��DJ�@�k{?1��e�[^_�Ð��������PS��  ������������������  ��������h\=�  ��������   �ƿb=�   ����   ��������hv�e  ������t`V�uh�OP�M�����Hu�E�     �@    �S������5��hR=Sh�;h�:�`  [^P������S�������&  ��E�    @�@�MXA룉�Q�u�uP�  ����t
�   ��������5��hR=Sh <떃�������hv�  ��XZ������h�H�  ���ۉ�tP��tLP�uh�OS�q�����H�5���W�uh�OV�X�����H�z������5��hR=Sh`<�������������hi=�!  ���������8lu�xlu
�x �����5��hR=h�<h�:�3  ZYP������S����XS������5��hR=hn=�΍v U��WVS��j 1ۋ}�k  ��;��}(1���������40W�G  ����uC�� ;��|�1��e�[^_�Ë���T3�L3�E��H�T3�E�L3�H��   �ːU��S���]j ��  ����x;��}�������]���1���U��WVS��j 1ۋ}�  ��;��}(1���������40W�   ����uC�� ;��|�1��e�[^_�Ë���T3�L3�E��H�T3�L3�E��H�T3�E�L3�H��   뻐U��S���]j �+  ����x;��}������D�]��Ív 1���U��WVS���u����}�E�t���u1��}� u
�? u�   ��[^_����������E��FG9�u����E�tŊ����u��1��ɐU��WVS���]Sh�=�u�u�}������1�Ht�e�[^��_�É����������u1���PWh�=V������H��   P�uh�=V�m�����H��   Q�E�Ph�=V�S�����Hu��E���������tc���������E��@u4���ًE�     �@    �    �G    �����1������K�������������E���������������������<����E� ��������t�����������������������������������'���������E�����������x���U��S���]�Y  ��Ph�=S�����؋]��Ív U��E� �E�E� �E�釮  �v U��WVS���
  �=����x�   �e�[^_�Ð��������P���    ���    �u���[^hzz������P�R���������$�����  ������ǅ���    ƅ(��� ǅ ���   S��$���h   W�>  ������  ��W�:�  ����������tm<#ti����(���P������P�����P��x���Ph�=W�O����� ��t[V�� ���h�=W��������������(��� u��(�����WS��  ���� ����U�����h8O��(���S��  ���ϡ�������� P�5�������ƣ�������x����$��蜫  ����������$�5�����|�  �D��������P�$�PR��P��(���P������P������ ��t����?�������������PR�PR��P������P��(���P�G����� ��u�������v ���������   ���������   h�=h�:�/  ^ZP������P�������(���PtUSh�Hh�:�  ��Ph�<h�:��  ZYPW�M����E�� ��u��W�������1��_�����W�����v ��6�h�:�v���h�j �5���5���+���� �����������P�'�����������Ph =h�:�j  ZYP������S�����}����u	��S�m�����S�w������U����ȍ��uUQjHh ��u�ȍ    ��  �������t
�   �Ív PjHh �hh����   ���  ���Սv �#  Ph>h�6h ��r   ����t���P��h�=h�:�
  ��P�\���U���hH=h>h�6�u�/   ����u�   �Ã�P��h>h�:�W
  ��P������U��VS��  jH�uV蚾  ���u�u�u�  ������tXPj VS�vx  �Ɖ$�\�������t9SVh+>h�:��	  ZYP������S�E����4$�����$�m�  �e�[^�É�1����h�@h�:�	  ��P��U��S���u�u�]S�������1҅�t ���t<
t�v C���t<
u�� �   �Ћ]��Ð�U���h�>�\�  �Ð�U��S�Ā�u��S  ���    �	  �}
  �$���  ����t4Hu�   1��]���PSh?h�:��  ZYP�]�S�T����$����PSh?�ٍv U����U   1��ÐU����܍��t�   �Ã�h�>h�:�  ZYP�5���J����$   �����$����������U������������    ���    � ����(  9�~����    ���    ���    ���    ���    �(  �d�   �`�   ��������  ��j�܍   ����1��Ð��U����!   ��t�Ã�h@?h�:�  ��P�l���U��VS��   ����t�e�[^�Ð��hzzhj?�P  ������t%P������Vh�=S�"�����Ht��S�?Q  ����뱃�V�إ  �����ڐ�U��VS��0�E�E���]��E�E ���]��]����E0�E��E8�E(���e������e����]����U����e@�������������������������ހ�E��@�UH�uL�MP�]T��   �E����e����������������������������������������
�E���
�E���������������1����]�uB����������u1�������������u��������u�   �ȃ�0[^�������������������E��������E�������������������E��@�.  �������������������ـ�E��@�
  �E��E���������E��   �}�f�E��f�E��m��]��m��E�P�$���]���]��E���������E��   �}�f�E��f�E��m��]��m��E�P�$���]��E��E���������Etp�E�����������Eu�ؐ������ ����E��E��������ـ�E��@u����E���   ��������E������ـ�E��@u�E��������ظ   ����������t��������6����v ����������������w������U���j�S�����1҅�t�     �@    �@    �@    ���ÐU��WVS���]�۸   ��   �E1��9�}%�P�U������M��4��u��������tF9�|�9���   �M1���t�}������1���эy��E�X����uN��~A���GP�����M���A������u
1��e�[^_�Ã��u�4���������   ����    ����P�h����U���Z랋}�W9��)  ����   �M�<�    ����AW�q�[����U�BXYW�r�J����M�A�}������}���   �E�X��tV��    �U1�������������Q������U��M���A�������������u�4�������}���������W�����U���Z�B    ��u�E�@    �     �������S�e����}�G    ���ӋM�Y�ǃ��G   j �-����G�$    �����G�����U�R�M�U��Y������U��WVS���E1ۋ89�}�p����4��u��������tC9�|�1��e�[^_�ËU�B��1��: ��H!����U��VS�u1�;|2���v����X�v�����    �F    �4$�����e�[1�^�Ã��F�4��n���X�F�4�C�a�����;|��U��VS���u�    h�q�u����������t=���uP���  ����t�����1��> ���e�[^�Ð��S������@u��ٍv �������U��WVS���}�    hzz�u�-���������t,��P���  �Ɖ$�A�������t
���e�[^_���������1�������搐U����U�<.t��u)��h�?h�:�   ZYP�5���I���������É�</t<"t<'t< ~<~B���u�   ��R��Ph @뱐�U����=`� t	�`��É���h�>��������t�8 u��6�܃�Ph`��*���XZhU@h`��	���붍v U��SS�`��ɋ]tJ��Sh`��d�������uQj�uS������]��Ã�Sh`�������Y���ZYPS��������΍v ��h�6j �����XZh�6j�����`�   ���U��S��  �Y   ��j P��� �������u�؋]���PSh`@h�:�=���ZYP��h���S�����$�������U���h�@��  �É�U��WVS��������E����  1���Ɖǹ��������щM�}�������у�M�Q������u�Vh�@P��� ����e��[^_�Ð�U��S��t�   ������   �����ta���    ��Shd������$d���  ����w
�d��]���Shd�h?h�:�F���ZYP�]�S�����$���������Shd���������u�봃�h�@h�:������P�ʐU���h�@�<�  �Ð�U��WVS��  �]�; u
1��e�[^_�Í�������A�   �ǉ������f�������� t�v �������������8 u������Ph�6h�6������V���  ���> t	�v F�> u�N�F</t�/F� ��������</t��uN��� j ���������������uX��j ���������������u-��j ��������������uB���t�CF뢸   ������������P�m�����뿃�h�  �������U�������������uh�@h�:����ZYPW������<$�W����v U��S��d  �uh�6h�6������S��  ��������PSj�������������t�Ћ]����w���9�����t1����&���1�9��������֐U��SR�����]t��x;�|1��]��á��������   �ڐU��VS��0���    �%�����Ph@Ah�6�&  �����ƍ]�t?��PSh�=V�k�����Hu��S��������x݃�S�p   ���σ�V�����������t	�e�[1�^��������P���=   Y^ShH=�̽������tӃ�hH=��������x���hH=�   ��뭍v U�����@����P�5���������X�u膙  ������D���1�É���U���塄������    1��Ív ��U��������塄���������1��ÐU����    1��Ð��U��S��  �u������P�uh�A�uƅ���� ����1ۃ� ��t�؋]��À�����iu�������nu瀽���� u޻   �׉�U��WV�}�uS�]� � �����t�v <@tB���u�1�[^_�Ä�t�9Ӊ�t
�C�A9�u�� B����BA��u�1��> tЀ? t˸   �čv U��S��  j@�]S�w�������t PSh�=������S�Ϳ���$���  �]����uSh�A�ܐU��WVS���E�E�    9E�}X�]�߉ސ�U�E��< t0�}tl�}~R�}t?��h�Ah�:� �����P��������E��U������9U�|��e�[^�   _�Ã�jW��  �ϋE��u���jV�l  뻃�jS�  뮐U��S��  h�Ah�:����ZY������PS萿��YXh Bh�:�k���YZPS�f���XZh`Bh�:�Q���ZYPS�L����$������U����u8���   ����1�@��B��v����1���@��B��v���   �É�U��VS�M�ɋu�]�Et#��P貮  �؉]�u���e�[^��'�  �v RPSV�   �e�[^��U����E���M�UtH��~3��t ��h�Bh�:������P�o������ÉU�M��   ����uΉU�M��   �U�M��4   U��SP�����]t�ۋM~�ډ�������Ju�[[���r�����U��SP�����]t�ۋM~�ډ�������Ju�X[���>�����U�����VS�ut%���]~����������S���Iu�[^�������ԍv U����E���Ut7��~"��t��h�B�p���1��ÉU��   �v ��u߉U��   �v �U��?   �v U��SQ���ҋ]t!1Ҋ���8uB��v�   �]���1����p����؉�U��SP�����]t!1Ҋ���8uB��v�   �]���1����5����؍v U��SS���ɋ]t 1Ҋ���8uB��v�   Z[��1���������ٍv U��U�E�E�U��3����v U����uj �u�u������U����uj�u�u������U����uj�u�u�������U��WVS���u�FP�}��  �X��<$�ݬ  H��9�!��    )�E��������e�[^_�ÐV��W説  H��PSh C�����������֍v U��WVS���M��u�E9E��   ���u�i�  1ۃ�9ÉE��E�    }I��1��   �;]|G�EE9�}=��+E�U�����	ǉ�CN��׋M���U��E�A9��M�|��   �e�[^_��;]}�P�uS�u�����������	ǃ��RP�u�u�   1��Ǎv U��WVS���}W�]跫  1҃�9E��E�    }+� �   9�}�u�2����BI����E�E�C9E�|Սe�[^1�_�Ív U��WVS���}W1ۋu�U�  ��9ÉE��E�    }.�   �v 9�}������U�C��I����E�E�F9E�|ҍe�[^1�_��U��WVS���u�]1����  ��9Ɖ�}!�E�؍H�   ;U��FC����9�|�e�[^1�_�É���   ����ݐU��WVS��  �u�]�}��������   �F���v������e�[^��_�Ív P������W������PS��������t �������PW�	���������   ��������S������@�����t�����PS�u������S��  ����t��j S�۵������t%���u�9�����h�  S�k�����P袴������VS腷�����=����E���PWh�C�5��藴��������Q������V������PS���������t��WV�:�������uE������RWS�u�6�������������������P�U���WS�u������S���  ��j �c���VWh�C�p�����U���j��������P�u�u�Q����Ív U���j �u�u�u�6�����U��SPj���a�����P�u�u����������xPjj S�2������؋]���U��VS�u�]j��������PSV���������x�E�q�E�e�[^�鬲���e�[1�^�Ív U���j �u�u�u��������x�Ezz�E��s����v 1���U��VS�]�uj��������PSV�\���������x#Pjj S�x����Ev�]���e�[^�� ����e�[1�^�Ív U��VS�]�uj���K�����PSV����������x#Pj j S� ����E�C�]���e�[^��ȱ���e�[1�^�Ð��U��WVS���uV�}W�:   ������x蠮  �e��[^_�É�PVW��h Dh�:�s�����P�b�����U��WVS��l  �c�  P������P�u�u�\k  �����ǋu�]t5��t������e�[^��_�Ã�������S������V�w�  �����  P��(���PSV�Q�  ���������x���SV�g  ���������������x���������u��(���B�҉�������  �x�9�8���tE��P�4:  ZYP��8����&:  �$�u�u�u��h@Dh�:�h�����P�W����*�������<����|�9�t��PR�u�u��h�D��������u�������  ��������  ��������  ������ǅx���cellƅ|��� ǅ����   ������PSV��x���P�������������������������������   ~���������1����$hH�����\������������������������V��    ������jH�����(���R��P���N�  1����������v ����������5t�F�Ѥ  ������P�~ڋ���������������������4�    ������蕤  ��p�����   ������P������P�uǆt�����ǆ���������������%  ����������l�R�,�  ���  ��������[��������������4�    ��p��u��l���������  �������������  ǆ�����������ǃ�  �������  �{  ����������  �����O  ���������֙  XZ�����������#�����t����  X�������+  ��  �q  �  X�������
  ���������  ����t,���  ����   P��x�P��f�P��4�P�K  �������������������������    ��������������h���t������������ǀ�      ǁ�      ���  ǀ�  ����u�����������j����S���  ��8�P蟯������W��x�P���������  ���������  �<������������7����n���Qjx������P��4�P茼  ���g�������l��u�����ǅx���fcelfǅ|���l ǅ����   ǅ����   �g���ǅx���fcelfǅ|���l ǅ����   ǅ����   �;����������u�u��h Eh�:�������P�Z���WSV��h`E����SV�u�u��h�E�Y����v U���j�(��u�,�    ���cell��� �$��  �ÐU���j�(��u�,�    �$����cell��� �w  �ÐU���j�(��u�,�    ���cell��� �$��?  �ÐU��E���1��Ð�,�U����u �E@���(�~�=(�v
�(�   1����(�   ��U��U��x1Ʌ҉�x���҉�tA��v�   �É����   ��U����0���t9���d�j�,��u�`��$����fcelf���l �y  �Ív ��h�H��������t�d�   �`�   띉��d�   �`�   녉�U����0���t9���d�j�,��u�`��$����fcelf���l ��   �Ív ��h�H蓪������t�d�   �`�   띉��d�   �`�   녉�U��WVS���u�}��  Y��Xj@V�\���1ۃ���t_���  �X�����$��  �YZPS�©��������t!��V�����Z�7��������e��[^_�Ív ��V觅  �U��4$�ؐ�E���0�C����$臅  ��Ív U��WVS��8�]S�
���������  P�E�P�E�PS�0�������t��Sh�H����������e�[^��_��蛘  �Z�  ��h�  P�E��ͩ�������E��  �}��   ~2���u��'���_�u�����^�u�����[�u��Ш���$ F닍v ��h���7����E���E�U����    ��h��,���l�ǂ�   �������  �U��$蹜  ZYP�5t�������t����  �v  ��jHhh�����P谷  ���}��  �E���E�U����    �}�$�����9  ǂ��    �E����U�E������    �����l��  �;  �  ���  ������  �}�5  �E���E�U�������E܍�l��E؋U؋E쉂�  ��p��E����  �E䉃�  Ǉ�    蘇  ��h�  P�E������������y  =�   ~O���u��h����4$�$���Z�E����  �Q���X���  �E���X���  �9���X�u�������$�H�������U䉗$�P��x��Ц���E؉}ԋ}�ǀ�      1���������Uԍ>���   F跛  ������P�~܋E���E�U���4�    ������ǆt�������p��t�  ��   �������u���������ua�E���E�U����    ������P��L  �������u�E����ǃ4�    �U�����������P�BM  ���у�����P蒣  ��닃�h@F����X�u�����X�U����  �ܽ��_���  �н��^���  �Ľ��Y�u������C�����h�Fh�:�������P��������  ����tDHt*P���������u����  ����������{��������P���������u��p�  �ԋ����$�������P�u��j�  ���7�������x�P�3  ��������j��t����   @P��p��a������  Z���   Y��   RP�e�  X�u�蘽  ��ǆ�      �|������  ���9�����j���   @P�
�����p����  _Z���   ��   RP��  ^�u��;�  ǃ�      [�u��x   �E�ǀ�     �$   ��   �j  �  ������h�F�K���X�u�����X�u�����X�u����������v ��S��h Gh�:������P�i����U��SR�E������������\�������t7�����u-���9�~$��~'��S�5���I������������v 1��]��Ã�S谺���݉�U��SQ�E@�t��X���9�~!��~$��S�5���������������1��]��Ã�S�_������U��SS�t�C���9�~!��~'��S�5��謺����������1��]��Ív ��S�����ݐU��SP�t���   ���9�~!��~&��S�5���[�����������1��]��É���S�ù���ސU��SP�t���   ���9�~!��~&��S�5��������������1��]��É���S�s����ސU����U�B����0�   w!1�������   �`��d��   �Ã�h@G�����������U��WVS��  �]S�uV�c�  ����u0PSV��h�Hh�:�������P�ʾ��������e�[^��_�Ív SVh�H������W���  YXj W�G��������   t�SVh�HW�ڶ  XZj W�$���1҃������U��WVS��  �]S�uV�Ƿ  ����u,PSV��h�Hh�:�?�����P�.���������e�[^_�ÐSVh�H������W�e�  YXj W诡������u��SV�*   ��SVh�HW�;�  XZj W腡������������롉�U��WVS��  �uh�H��x���S�����uhIS������S��  ��j S�4�������t-��S��hIh�:�s�����P�b���������e�[^_�Ð����t���PS�$�����p�����t�������t��S��hI뮍v ����p���h'Z�����������l�����   ��P�_~  �1I��l����   ��������8¾   t"��l����8I�   ������8¾   ul����p���h>I�U���������t;��P��}  ���;xu�{du�{ru�{ t�P��l����uh�G�X���������p����W����������PS��l�����h�Gh�:�.�����P����X��p����!�����������v U��VS���]�uS�0�������x0��u�]�e�[^������v ��V�s����$�+������e�[^�Ã�ShII�w����v U��VS���]�uS���������x/��u�]�e�[^��+����v ��V�����]���e�[^��R�����S��hIIh�:�P�����P�����v U��WVS���}�������������t��h H����������e�[^_�Ã���x�V�Q,  �E� ������   �U�B �@�Rl�\��9�r'�P�s�s�s�s�s�3V�T1  ���E�� ;Xls�Q�u�V�]�S�u�e0  ����~#�����u���u���u���x�P��/  ��RVS�u��0  ����~#�����u���u���u���x�P�A0  ��1��'�����V��+  ��U���8�    1��Ív U�@����VSuu� ���jV�]�  �H��@������5,�u1�����jS�5�  �s�    ����H��e�[��^�Ív ��j足���Ã�����X뻍v ��j蚳���ƃ��,��p�t���U��VS�<�����   �@���j8S蹍  �H��C    �C    ���<����C    �C$    �C     �C0    �C    �C    �C,    �x�u1�����jV�Q�  ��F    �5���H��e���[^�Ív ��j�Ҳ���ƃ�����p뻍v ��j8趲���Ã��x��X(�4���U���jh|���  �|��Ív U��WVS���E��E�    1��E�    �E�   �D�����������щ˃�x���</��  Ky�@���t'���N��t�F$��t
�8����  �F�F �v(��uۃ}�}  �M�Y�޿3M�   ����   �޿2M�   ���   �޿1M�   ���   �޿8M�   ���  �MtT�E�E��;-��   ��j=S�  ������   �E���t�=<�����   ��j=S��  ����tK�Mu��w  �  �}�E��t(��  E�u��u1��v �e�[^_���  ��������  E���VSh�Ih�:�����ZYP�5��菙���E�   ��늃�S�bu  �\��E�    ���S�s  E���C����Z����v ����P��  E�C�����u��9����Y  �i����8���u'�}�p�����j �+������������7����v ��j ��������tȃ��E�0�n  ���E�   ������v �1����������Q�����FXZ�F$�0�v�����V$�B�����   ������v �~�1��������ы<��M�������у�M�Q�v�/����FY_h8OP蛚��XZ�F$�4��v苚��C�V$������u��l����T�D��:����U��WVS��  �D�����  �|����D  ��hPMh�:�,���Y[P�5���җ��XZj�5D���
  �������@�����td� ���ƅ���� ƅ����[ƅ����-�   t�����*�����B��u��Ƅ����]Ƅ���� ������������P�j
  ���������<���ǅ����    ��   �@�����   ��C����u�{�]  �<b1��;��������эQ�;�����~������fǅ����  �C���	  ���3������P����Y_hZM������P�	���XZV������P������C������  �C���a  ��������������P�	  �[(���ۉ������@������5��j
�X����@�������   �<���u
�e�[^1�_�Ã�h\Mh�:�n���ZYP�5���@���������tʃ��s�3������hjM�5�������C�� ��uD�C ��u	�[(��u�뒃�Phd������hvMh�:�����^_P�5��褕���� �ƍv ��P�������Q  ��먃�h�Mh�:�����^_P�5��� ��c������������w�Ph�M�5���A��������u����������h$n������P�l�����������h�M������P�P���Y_V������P�A���XZh�M������P�.������:�������h�M������P�������������d������h�Mh�:�����^_P�5��莔�����5|�h�O�5���u������{����P  ���D��\����D��M�M���U��VS�]����ut,�v �Ѓ�<tP��<7��&t��V��P����C�����u׍e�[^��Vjjh�M蹗���ލv ��>u�Vjjh�M��v Vjjh�M��U��WVS��,�D����]  �5��j'jh�I�i����5��j-jh J�U������5D�h�M�5���|����|�������  �<�����   �E�@��Eԅ���   �UԋB���8It����  ��MHt�0]�Eԃ��x�Z  ��MP�Eԃx�;  ��MPR�U��2h@J�5�������Eԋ@�� ����  �Eԋp����  �UԋJ,���  �Uԋz ����  �UԋJ����   �Eԋ@(�5��jjh�M�E��A����Eԃ����'����=@���tF� ���t=V�Ph�M�5���K����K����u=�[�5��j	jhN��������u��5��jjhN�ϕ���e�[^1�_�Ð�5��jjhN谕��XZ�s�5�������5��jjh3N茕���� 농v �5��jjhFN�p���XZj�Eԋx�1���������Q�$���^�ǋU�X�rW����Y[h8OW����������tP���5��j
jhRN����XZS�5��������5��j	jh]N�������h8Oj 跔��������u��5��jjhgN�ʔ���<$�������\������5��jjhtN褔��[^�E��p �5�������5��jjh�N�}����� �	������j�EؕN�EܙN�E�N�E�    �z,�1���������Q������XZ�E��p,W�Δ��[^h8OW�����5��jj��h�N����1��� ��t�M؅�u'�5��jjh�N�����<$�;������]����v S�t��h�N�5�������XZh8Oj 聓��F������t��D�؅�u�뢐�5��jjh�N舓��Y[j�Uԋz�1���������Q�<�����XZ�E��pW�����[^h8OW���������þ   tN�QVh�N�5���n���XZS�5�������5��jjh�N������h8Oj �͒��F������u��5��jjh�N�ߒ���<$�3������G����v �5��jjhN踒��_X�U��r�5�������5��jjh3N葒���� ��������N���������N�������0]���v����5��jjh O�O���XZ�5|��5���0����5��jjhO�(����� ������C  ���D�������D��M�����v U��WVS��$  �u������S�u�~���hdVh$Oh�:�U���ZYP�5����������� �������������������v ��j,���������  ������tv� 1����������������Ӌ��������L*W������h6O�5��F芍���������������뙐hd������Qh:O�5���������V������1���������������ы������L���L!V������h�O�5�������e�[^1�_��hd������h:O�5��������뿍v U��WVS���u��1��������U�хҍy�~�ύ:��L~��u�����5��V�i����e��[^_�Ív �5��jjh@O�H������ɍv U����@����Mt9� ���t��9�t �R��u�PQh�J�5���D����   ��1��B��PQh�Jh�:�p���ZYP�Ѝv U��US����]t��9ع   t	B���u�1ɉ�[�É�U��WVS��\�u�<=�U�t�v �F�B<=u�� 1��E�    �}���������ѻ@�IF�ۉM�t>�v P�u��3�E�P腍������u�E�1��]��;���������I;M���   �[(��uŃ}���   �E���t}�U��B4@�B4Ht_�z1���й�����ˉ����������у��Q�E��p�����U��BY[h8O�r�W���XZV�M��q�I�����1��e�[^_�Ã�V��f  �U��B��P�M�Qh�Jh�:����^_P�5��蹊���   �P�U�RhDO���E�   �1�����U��WVS���<�1���u1��e�[^_�É��@���t1�v �C��t�C��t�s��tQ�C$�1���u$�C0��u�[(��u҉�븉����s��ǃ����4��s�s�3�(   �F�C$������u��P�s�s�3�   ǃ�륐U��WVS���E1ۃ��}�u��   ����   H��   ��tj��~
��t4��t
�e��[^_��VWh Kh�:�����ZYP�5��膉�����ҐWVh@Kh�:����_ZP�5���a������uh_O�PWh�Kh�:����Y^P�5���5������uhwO늃��uV�4   �Ã��O��������D������uV�W  �ݐ���uV�  �Ή�U��VS���E�Ph�s�u�]�̋����H�   t	�e�[��^�Ã�j-S��������t8�E�P�E�Ph�OS蓋�������   uŋE�;E�|	;E�1�봺   뭃�j,S�G�������tL�u�PVh�sS�L�����Hu)�E�9E�tŊ��t�<,tC���t�<,u���t�C�; u�먺   �R����v P�E�Ph�sS� �����H�   �0����E�1�9E����������v U��VS��$�E�Ph�O�u�]�������H�   t	�e�[��^�Ã�j-S��������tL�E�P�E�Ph�OS臊�������   u��E��E�������Et�E���������Et1�뤺   �������j,S�'�������tX�u�PVh�OS�,�����Hu5�E��E���������E��@t����t�<,tC���t�<,u���t�C�; u�똺   �2����v P�E�Ph�OS�ԉ����H�   �����E��E���������E��@�������������U��WVS���]�; �uu1��e�[^_�É���j,S�]�������tq1������������PIQSV�J�������u'1�����������р|�,t����������р|� t����t<,t��C���t<,u���tC�; u��   �s�����SV�ǅ�������������W����U�<���V1���Su1��e�[^�Ív �@���t�v �C��t�C��t�[(��u���эv �s�3h�Kh�:�����ZYP�5���~���F����U��WVS���<���t%�E�@��E���t�E��@��u�M��I(�ɉM�u�e�[^1�_�Ã�j(�E�
   肜���U��z�B$�E�    �     ���E���1�����t<,t��C�F��t<,u���FP�<������M�U��VW�M��A$�U��4���  �M��U�A$��� B�M��9ʉU�}.�M��A$�U�E���    �; �9����{ �{�r����'�����
�ȃ���P�E��p$�M��/����U��B$���U��WVS���<���u
1��e�[^_�þ@�1���tP�N��tB�F��t;� ���   t�<,��   B���u�F$�1ۅ�t
��C����u��ؙ����u�v(��u����Q�6h Lh�:����ZYP�5��贃����Sh@Lh�:�����ZYP�5��蓃�����vh�t�5���}���G��똍v A�j�����U��SP�H���t9�����C��u!���t��P�   �[����u�1��]��Ð��P�#   ���5��j&jh`L�ц���$���������U��VS��  h�Lh�:�u�3���Y[P�5���ق�����v������h�OS�r���XZj S�s  �F�e�[1�^��U��WVS��   �u�vh�Oh�:�׿��ZYP�5���}������6h�Oh�:赿��[_P�5���[����F������  �F ����  W�^����  ��OPh�Oh�:�m���ZYP�5�������F�����S  �F���!  ǅ����    ��������ƅ���� �^,����  ��WV�  ������������   �F��tWP�v�6���������Q  �F0��t��W�Ѓ�����   W�6h�O������S�!����F,������   PSh�Oh�:螾��ZYP�5���D���YXj��h�Oh�:�z�����P��q  ����uj��������u4�V��t
��������tE��u��������~�V��u&��u
�F��t�v ������������F��������e�[^1�_�Ã�j�蔃����S�������������PWhPh�:�۽��Y[P�5��聀��Xƅ���� Zj��h!Ph�:谽����P�'q  �����h���됉����ύv ��h0Ph�:�~���ZYP�5���$������5��h   W���������t&����������������<
tB���u������ ���j� ���QPh@Ph�:����_ZP�5�����������Ph�OhNPh�:����[_P�5������������\P�L���SPh}Mh�:踼��ZYP�5���^��������QPh_Ph�:葼��_ZP�5���7����������v U��WVS���   �M�Y,����U�t�<,t
�C�B��u�� C�����h���t��<,t
�C�B��u�� C�����(���t��<,t
�C�B��u�� �A���T  �]���ou�}�lu�}�du�}� ��   ����nu�}�eu�}�wu�}� ��   ���H�}��   ����   ��au�}�nu�}�yu	�}� t9�v S�E�Ph�L�5���3~���5��j0jh M�߁��������e�[^_�Ã�j��(���P��h���P�uh�6�s  �Ã� ��t1��ˋE�  ��(���P��h���P�uh�6��s  �Ã��΍�(���P��h���P�uh�6��r  �܍�(���P��h���P�uh�6��r  ������t���P�u�"���^_P�u�Á��롐��hmPh�:蚺����P�s  �������U�����    �ÐU��WS�]1�����������эy��������9�}0��S��R�P�������������� �e�[_�É�����   P�5�����艔����������륐U��WVS���E�E��E�    �E�    �1��ۉ���   �E����   �M�|��������9���   ����'����u����t"��'tS����������F�����uދE��t�������'���������� �e�[^_�Ív �������'\''�D ���롃���   ���P�5���y������������B����E��E�e�[^_��T�������E�M��Ӌf�P��f��u��Rh�P�z������t��'tF�G��u��������E����E�   �߉�U��VS��������  �$������@�����t� ���t��{ ��   �[��u�<���t�@���t��s��u�[(��u򡐵�e�[^�É���hd����Y�3�{����$ZM�o���Z�C$�0������C$�@�����   t�����h8O�C���X�C$�4�����F�C$������u�낍v ���hL��N��������B���U��WVS���u���}�M~v��~r������    �Й���Å�~9�}
T�9�~PSh�P�5���T���y������c�e�[^1�_�É����5��j
�{���T��������Ր�d   뛐U��WVS���5���}��y��Y�5���u���y���4$�z����1҅�x;�<rtG�]�<rt8�u��dy����t91҃��t��V�����y��XZWS�x���e�[^��_�Ëv�ƍv �]�뷃�S��x��1��?r���$��x���4$�v|���4$��x���$    �uh QhQhQ��w����j�|����U��WVS��(�]S�rx���ǉ$�H{��^Xjj��x��Y[jj�E���x���E�XZjj��x���]�E���މ���S�u��|����;�����t:@u��E��������u�j�x��_X�u�j�wx��[^�u�j�kx���E�e�[^_��@u��Đ��U��`��É�U��WP�U1�����������щȃ�x�v �</tHy���R��S  �`��}�1��ÍT��U��E���dP�8  �E���U��U���   t��~���   t�   ��t�������1������U��E���UtJ��~1��t��t1��Ív �Ҹ�Qu�Q��Ҹ�Qu⸴Q�ۅ�uՅҸ�Quθ�Q�ǅҸ�Qu���Q�U����U����Qt���Ҹ�Qt
J��Qt1��Ív ��t��cu��h�Qh�:�����݃�h�Q��U��SP�]�������vVh   ��h����Qu��QPh@R��  ����u���۸�Qu��QPh����z��������]��Ív ��SP�����$�������U����m�����w��P�����Ðh   h��h�dhR=�_  ����t����֐��hKRh�:�6���ZYPh���=z������U��VS��  h   ������Sh�Q��h@Rݝ������   ����us݅������������t
�e�[^�Ív �؃�j ������ơ������t%1ۃ�����V��   ����u��������u�݅�����݃��ݕ����롍v P������Ph�OS�x�����r����U���h   h��hcRhR=�I   ��������H%���É�U���h   h��h\=hR=�   ��������H%���É�U��S��  hH=�uh�6������S�%�  �u�u�uS�ƞ  �� H�����]��Ív U��WVS���}���ut]��tY���t	�> u��u�> t1��e�[^_�Ív �   ����P�0   ����$�#   GF��9�uɊ��t��> u�볐1�9���봍v U��U�B�<w�� ���Ð��U��E�@     �@    �@    �Ív U��S���]S������K����~���sl�v�����S|��u�C    �]��Ð���sp�}v��X�st�tv���Cx    �C|    ���̐U��WVS���}�W ���   �����	�Ҹ����u�e�[^_�Ã�jQ襊���GpXZj�G ��P蓊���Gt�G ������  �Wl�@�\��1�9ӉU�rA�Op���h  ��A��������ـ�E��@�G  �F���C�S����QF��;]�swxh�,jV�wp�kt���Ox1��A���9���   �w����   �G<�W@���   �GL���   ���   �_��t0��t�GD�WH���   ���   �GP���   �G|   �   ������Gp�T�����D�����   ���   �E�jP������E����   ��뼅�t�Gp�P� ���   ���   ��j�E�P�Ʒ���E����   ���Ox�\������Gp�D������(7�$W�h  �Wt�Ox��F�A���9�|�������v �������������Ox������U����E�@|    �@    �     �@    P�^����   �Ív U��E� �É�U��E�@�ÐU��E�    ɸ   ÐU��E�@   ɸ   �U��M�E�U�AT�E�QX�U�A\�E�Ad�E �Q`�Ah��U��S���M�A ���E�E�]�E ��  ��������E�AT��  ��������E��  ���]��ʋE�U�AT������E�QX�A\�_  ������E�.  �������]�U�E�Q`�Qd�A\R�$�$�$����������E��   ����������E��   R�$�}�f�E��f�E���m��]��m��E��Qh�AdR�����$����EuS������Eu"����R�$���m��]��m��E��Ah��[�É�������Eu���m��]��m��܉����m��]��m��͍v ����뫉���������Eu���}�f�E��f�E��m��U��m��d����}�f�E��f�E��m��U��m����G����v �������������v ��������Eu�����]������������]��������������v ��������Eu���U����`�����U��W��������������:�����A�������A�����������}�f�E��f�E��m��] �m���[�������U��WVS���M�A ���}�]�u~0�AT�QX�W��A\�}�Q`��Ad��Ah��W�   �e�[^_�ËA��uɋA��u�jS����XZjV����Y[jW�s���XZj�u�g���������U��E�@ �ÐU��EVS�U�@�rl����L�]��K�T�L�]��K�U�L�
�T�E�[^�Ív U��SP�]�C9C |��u ���C2   h�  �Є���Cl���]��Ð��2�C�@����P�sl�$����ډ�U��SP�]�E�U�M�C<�S@�KLQ�$���$QRPRPS�a����C|�� ��t�C<�S@���   �CL���   ���   �C   �]���U��S�]�S��u
1��$�Ív �S<�E�K@�H��E�SL��   �ۍv U��SS�]�E�U�M�KP�CD�SHQ�$���$QRPRPS������K|�� ��t�CD�SH���   �CP���   ���   �C   �]���U��S�]�C��u
1��$�Ív �SD�E�KH�H��E�SP��   �ۍv U��WVS��(�]�E�E��S�]��]��}�u �Z����C �@�Sl�E��E��ɍ���������uf����Z�z�r�C|��u*V�$���$W�u��u��u��u�S������C �e�[^_�É����sp�n��X�st�n���C|    �Cx    ��믐�����E��E�����Z�r�z뎍v U��S��$�E�Xl�@ �@�L��9�ss���S�E؋C�U܋S�E��C�E�C�U�E��Q��A�S�Q�C�A�C�A�S�C�E؋U܉�E��Q�U�A�E�Q�A�E�A����9�r���$[��U��S���M�U9��E�E�E ��tP��������E��@��t8����)�R�}����$f�E��$��$f�E��m��]��m����]�؋]��Ív ����������������U���E�E��������u�   �Ð1���U���E�E��������Eu�   �Ð1���U��WVS��H�E��EP�U��]��}�f��������E���  �7��t&���}�f�Eڴf�E��E��m��]��mڋEԍe�[^_�Ë_��t5������������Eu�(7�}�f�Eڴf�E��m��]��m����%(7���G ����  �O|���`  �Op�������Eu.݇�   ������u	���   끐���E�jP�2����E��j����wx�D������������Eu݇�   ��������uŋ��   �:����V�����������E�    �űGt������   �<)���$�t��t��]��փ����E���   �Gp�t��4؃��$�]��փ����E�tK�ډ]�UЉ�������Op땋Gt����t$���$�p�p�p�p�p�0������ ����݇�   ������t݇�   ��������������������C�U�ډ]�덐�)�9�����W�]����������E�������G ��~$���$W�]��  �����E��]����������G��t�G<������u
�؋GL������G��t�GD������E�M����GP��������>������O��u�W��t%��������w��������_����������	�������������������U��WVS���E���u�}~.�Ã�V苮������u$P�v�6�u������������Kuԍe�[^_�Ã�jW���ެ����U��WVS���E���u�}~0�Ã�V��������u(����$�u�����������Kuҍe�[^_�É���jW���~�����U��S���]S������1҅�u'�E�� ������E�����t��������E��@���ЉЋ]��Ð�������U��U�B �Jl�@�T��9��Er6�������������u�B������t��9�s���9����!�����������U��VS���  ��(���S�u�^����$������S�uV��  ����x�   �e�[^�É�PVh�R������S�-i���$蹂��������Չ�U��VS���  ��(���S�u������$�N�����S�uV�  ����x�   �e�[^�É�RVh�R������S��h���$�Q���������Չ�U��WVS��p  ������V�u�}W�]  ������   S������P������SV�9  �$�5�������u��������P��������t(QWh S������S�=h���$�Ɂ��������e�[^_���u�u�������������������������uW�   �ύv VWh@S몍v U��WVS���  ������ESݝ����u�}�������u$�u WV����������S�������S�u�u�9   ����x�   �e�[^_�ÐW�uh�S������S�sg���$������������U��WVS��d  �uV�]S�}�p�������u5WSh�Sh�:�̠��ZYP������S�!g���$譀��������e�[^_�Ã�������P������P������P������PW������WVS�<�  ����x�   �VSh T닐U��WVS���]�}�uS�����]�u�}���e�[^_�� �  U��S���   �u��(���h�HS�vf��XZhfUS�"  1��]��É�U��S���]Sj��  YXSh�   ��  1��]��É�U��WVS��  �u�u�]�	  XZSV�=�������u^P�E�PSV��  ���������x�E���t�   �e�[^��_��P�u�E؃��$�  ���u�E܃��$�  �   �ɍv PVh�H�����P�e����ShfU�����P�������������uH��~��W�a����SVh@Th�:�����ZYP�����P�Le��X�����P��~��������K����WShfU�����P腭��������x�=�   ~ ��P�8a����hnUh�:蒞�����Qj������PW�Qe�������   �����jj������P��x���P�c��XZ��p���P��x���P�c��������������h���P��x���P��b�����������S�u��t�����p����;  ���u��l�����h����$  �<$�t`�������v U��WVS���  �u�]�  XZS�uǅ0���    �8���������  P��h���VS�u�0��������m  ��V��������u��V���������   P��H���WS�u�|���������   P��@���P��8���PW�X  �4$��������tmٽ6���f��6����݅8���f��4���٭4����]�٭6���݅@���٭4����]�٭6������u�u���  _X�u�u��  �   �e�[^��_�Ív ݅8�������������EuN�(7����ٽ6���f��6����f��4���٭4����]�٭6���݅@�����������Eu���j������c����(7��밐�����뀃��E�P�U�R��@���P��8���PV�V����� �9�����S�uh�T�����S�gb���$��{��뱐V�uh�H�����V�Gb����ShhUV�ȃ������u=��0�����t����0����	a����S�uh�Th�:蟛��Y[PV��a���4$두QShhUV����������0���t�RPh�   V��_�������   ��������E�P�E�P�E�P�U�Rh�UV�E�    �E�    �E�    �E�    ��`���� �����E���1�9�}$��~�D�؅�t���u�t����  ��C9�|܃���0����.`���   ����U��WVS���   �}����[^PW�?�������t\��h U�����V��`������hhUV�+  �қ��PWh@Uh�:�q���Y[PV��`����V�Wz��������e�[^_�É�QWh�H�����V�`��XZhhUV�L���������t��E�x��t��S�h_��1�붋E�p�0h�US�\��^����U��WVS��p  �uh�H�����W�<`��[^hfUW�o���������xG�E�H��t��S�C\��1��e�[^_�Ðj j������P������V�Q^��XZ�uV�V^������u?��hfUW�  踚��P�uh@Uh�:�U���ZYPW�_����W�;y�������돋E����PV� ^������t�Wj������PS�i[��^�Z����v U��S���EP�]譢������u�C��t�E�C    ��C1��]��Ð�E;}�;C���U��S�� �E�E��E��UP�U�]�Ѣ������u�C��t�E��U��C    ��S�C�S1��]����E��������Eu��C����������Eu�[�ԍv ����U���j �u�u�u�   1��É�U��WVS���]��K���u�}~F�v ����E��E�P跡��������u!�M��t>�E���t�W��t �G    ��G��K����e�[^1�_�Ív ;}�;G~��܍v �E��čv U��WVS���u����N���]�}�]�~N������   ����   ����   ��WS�Ǡ������u^�E�P��t"�E��@    ��X��N����e�[^1�_�É��E� �E���������Eu=�E��E�@�E���������Eu �E�X��W��M  ZYPS�  �Ã�뢐����������]��e��������[��������]��M�����U��S���]jS�b���YXj�CP�U����C   1��]��Ív U��WVS���]�K�ɋu�}t#��jV� ���XZjW�������e�[^1�_�Ð��S���������u(�����CP��������u	�C��ǉ���뵍v ��jV�Ş������U��S���]jS����XZ�CjP�	����C   1��]��Ív U��WVS���]�C���u�}t#��jV�Ԟ��Y[jW�ʞ�����e�[^1�_�Ð��S迟������u4��S�V����CP袟������u�C�S�W�뻉���멍v ��jV�m�������U��EE�ÐU��WVS���]S�uV�}胞������t ��SW�r�����������J�e�[^��_�Ã�SW�R��������   u���tO��~2��t1�������������Eu���غ   �������E��@��렅�uϋ�9��   �9��������������Et����������뷍v U��S���u�]�:K  �؃�S�u�u�Tf  1��]��ÐU��WVS���E��uP�}�]�u��ޝ������u;��t*��~��t�e�[^1�_�É�V�$����鐅�u�7��V�$����ՐPSjW�.�����U��VS��,�E��EP�U��]؋u�]謝�������E�uB��t9��~��t�؍e�[1�^������t�����}�f�E�f�E��m���m��Ԑ�����RSjV贛������U��VS��<�E��EP�U��]ȋu�]�l��������E�uB��t9��~��t��1��e�[^������t�����}�f�E�f�E��m���m��Ԑ�����QSjV�8��������뾐U��VS���]S�uV�+�������u\��t;��~.��t	1��e�[^����}�f�E�f�E��m��]��m�E��܍v ��uӋ����}�f�E�f�E��m��]��m��։����E�jP�����E�뢐U��VS���]S�uV蟛������u0��t'��~��t	��e�[^����]��E������u��������j�E�P�����E��ΐU��VS���]S�uV�?�������u(��t��~��t	��e�[^�������u��������j�E�P����E��֐U��WVS���  �E�     �@    �@    �@�����@�����@�����@    �@    �@     �@$    �@(    �@,    �@0    �@4    �@8    �@<    �@@    �@D    j j �uǅ@���    �.U����ǅD���   �R�uh   ������P�+��������0  ��@��������  Q��H���P�����S������P�  ����tI����   �޿i=�   ��u{��@���   uL�E����P��H���P�1  ����t��@�����D����X�������D���������P�C  �e�[^_�Ã���D�����h�Uh�:�������ҍv �޿�y�   ��u���@���   u)�E����P��H���P�  ����t���@����o�������D�����hV땍v @�����X�����@���   ��  ��@���   u��j ��h/V�X���Pj j �u�S����ǅD���   R�uh   ������P蓅��������  P��H���P�����S������P�  ����tn���V  �޿i=�   ��tU�޿�y�   �tE�޿BV�   �uY��@���   u4P�E�p��(P��H���P�n:  �����g�����@�����D����E�������D�����hGV�m����v �޿]V�   ��uO��@���   u+P�E�p��0P��H���P�:  �����������@���딃���D�����hbV�������޿xV�   ��uS��@���    u.P�E�p��8P��H���P�,:  �����������@��� �1�������D�����h}V�����v �޿�V�   ��uS��@���@   u.P�E�p��@P��H���P��9  �����9�����@���@���������D�����h�V�E����v �޿�V�   ��ug��@��� xFW�E�p��P��H���P�C:  ����������E�@���������������@����   �T�������D�����h�U��������޿�V�   ��uk��@���   uFV�E�p�� P��H���P��9  �����]����E�@ ���������H�����@���   ���������D�����h�U�Q����v �޿�V�   ��uc��@���   u>�E����P��H���P�  ����������E�X���������@���   �e�������D�����h�V������v �޿�V�   ��uc��@���   u>�E����P��H���P�  �����n����E�H���`�����@���   ���������D�����h�V�i����v �޿�V�   ��uO��@���   u,���u��H���P�!  �����������@���   ��������D�����h�V������޿W�   ���������@���   u0�E����P��H���P�  �����������@���   �'�������D�����hW�����@������d�����@���   ��   ��@���   ��   ��@���@   ��   ��@���    ty��@����  t[��@���   u��j ��h&W�,���P��@���%   P��@���   ��@����u�>  ����t
��j �����1��������j ��h9W�������j ��hLW�������j ��h_W������j ��hrW������j ��h�W������j ��h�W�����U��WVS���]Sh�`�uV�}�.O����1�Ht
�e�[^��_�À;#t3WSh�WV�
O�����������u׃�S�*  �<$�*  �   뿐1��U��S���E�P�uh�W�u�E� ��N��1ۃ�Ht	�؋]��É��}� u�   ��v U��S��  �E���Ut0RPh�Wh�:�ǈ��ZYP������S�O���$�L'  �]��Ív SRh�W�ې��U��WVS��(j �}�E��  ��h���E�M������  ���E�P�E�P�E�P�E�P�u�"  �� ����  �u��u��u��u��  �ËE���9E��  ���M  ��h�]  �$b���U�������   1��E�    �E��]  ��S�u��  ������   ;u���   �M��uF��G@����������t���Ív �G8������u��C�G(������t����G0��������u��U�
�C8�U�ЋE��\���C�\���E܃E�F�b��������u؋U�2���  �E���a���U������W�����h�Xh�:������P��f�����u�YL���$   �Ag���U����u
�e�[��^_��Pjjj�Y���������5��j
�xK����h�Wh�:貆����P�f���������E��@P��h@X�i�����h�X�\����v ��h�Xh�:�j���[^P�5���I���������U��VS���u�u�  �Ã��۸����t*P�u�uS�>  �Ɖ$�pK�����������x1������e�[^�É�U��WVS��$  �u������P��L����j@������R��G���� ��t�  ��������P�u��襆����Ph�X������S�L����hzzS�K���ƃ����������  �E��t	�U�    ǅ����    ����V�oG���������  WVh�   ������R�I��������   ������1����������I1�1�9�}9���*����<#t-< ��   <	��   <
��   < t<	t��=����GB9�|ȅ��p���Ƅ/���� �E���������W�������������S�E�0�,_���U�؉������G�$�^�����������B�W������P�U���p��}J���E�C�� �����������[����s����]��t�������E���������t4�U��t-����������������S�E�0�^���U��D�    ���������e�[^_�ÐU��WVS��   �}W�u�]�  �ƃ��������t0P�C2PSV��   �����Cd~zHtf�������V��H������x�؍e�[^_�Ív ���t4W�uh Yh�:�l���ZYP��x���S��I���$�Mc����������W�uh@Y�ʃ�SV�  �Ã�뎃�V�zH���Cd뒐U��SP�]�{dt
1��]��Ív �Ch��~���st��]�����Ch    �؉�U��WVS��  �uh�   ��h���P�,G����1Ʌ���   �   ��h�����Y������1�8���   �E�  �E�  ǅd���    P�uh�   ��h���P��F��������   ��h���P������Sh�Y��h���P��G������uk�޿�Y�   ��tb�޿�d�   ��uI����h���P�u�I����d�������d����o����E�8 t�E�8 t�   �e�[^��_�É�������퐃���h���P�u뭐U����u�uh�Y������U��WVS��  �E�xd��  �@p�U9Bl��  �Bh����  ���u�  �������E  Pjjh�Y�G�����uh�YW��C���E����2Ph�YW��������C���U1��Bh��9���  ��Kx���U�Bt����P袊������tKy�9��4  Wjjh�Y�AG������W�F��Y[�u������V��G����j@V�B���� ��t�  ��V���������y�����Ph�X������S��F����h�YS�F���ǃ����   ��   Rj j W�}D��蔁��P�uh�YV�F���� ǅ����    ��W�3B������u5PWh�   ������S�iD������t��SV�xB������u�ǅ����   ��������t��W�$E���   �e�[^_������P�uh�YW�cB�����щ�P�U�Bl�Ph�YW�GB�����U�Bt����P�2�������tP�5��h�OWF�B����9�~�����P�U�Bt�4�h�U�܍v �U�Bt����P��������t�UF�Bh9�|������U�Bh�	������X�����P�u��h�Yh�:��~����P��^�������������h�Y���hZh�:��~����P�{^���v U����uh�Y轍���Ív U��WVS��   �E�@l    �@t    �=��������1����I1���h�����\���ǅ`���   P�uh�   V�B��������   ��`�������   Q��d���Sh,ZVǅ`���    ��C����Ht{R��\����5��V�B������u?��jS蜆����G����    S�E�pt�RX���U�Bt��d����T����^�����PSh�sV�WC����H�����t��e�[^��_�Ë�d����U�Bl�)�����d����i����U�Bl�H�Bp�zh�   ��U��WVS��x  �]S�|�����������xb�~��Q������V�Ǎ�����PS��������t��VW�?�����������u)��j RWS�u������S�;U  ��P�@����1҅�t�e�[^��_�Ív ��S�@�������   tރ�j'S�>�����������u�PSh`Z������S��B���$�Y  1҃����T�뜐U����u.  PjHhh��u�]N  �   �É�U��WVS��j j �uV�0  ����t��Ph�Z�\��������e�[^_�Ë=���������~���1�1ҍv ������   C��(  ���   ~��~ ��Q�A  ����������������RjHVhh��M  1����   ����������tU��tP��tK��tFC��(  ���   ~��z:  �����d���诛����j蹚���$   譚���   �����v �>u���S�)  ��말�F9� �t#9��&�����h�Zh�:�{����P������F9���u��������U��SS�]�K��u=�S,��u&�C4��u��S�U���]��Ð���s8�U��������s0�qU�����ʃ��s�aU�����U��WVS���}�p  �E���e  �E���Z  ��j<�iT���ƃ�1�����   �E�F�}�    �F$    �F(    �F �F    ��   �E���F�E��~�E����P�T�������F8��   �E�F4�E��~ �E����P��S�������F0tN1�;}|�U�V,���e�[^_�Ív ���^0h   �S��������tG;}|���OuG���v0�PT������}��~���v8�:T�����}��V�(T��1�뙃��v�T��������F0�4��T����Ou�룉��U��������P�)S�������F�����먃�h [��X��U����������P�u�u�   ��U��WVS��@  �u������h   Vǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ��<���������������tF���#t�6?��� ��f�P%   f��u1��-t,��+t'R�uh   W�<��������u�������e�[^��_�ú����1��������р|�
��  ������S��h���Wh�\V�=����H~,P�E�u��PS�#  ����tP�u�uW�$  ����uSWh�\�5���j:��������t�����j|V�}a  ����������Y�����j|�@P�_a  �����ƺ�����9���F�> �  �������U;B���  P�B��������Ph�\BV��������<������������������j|V��`  ������u������ty�Ѓ�%��  ��%�.  ��#��   �������E;P,}5��V��  ������~;PSV�U�B0�������4�B���������  ����V�i  ������t���u��E�x�t
��������t1�������E;P|#������;P,|������;P4|�������������������������u�U�B��tZ��~A��tǅ����   �o����ES��$Ph�\V�;����H�R���ǅ����   �C������u�P�E��Ph,Z�͐�EW�� Ph�\뽐��@�������t�~ tF������U�z�t���������J����������U;B�8���������;B,�)���������;B4������������E;P4|"ǅ����   ��V�  ������������F�������8���U�     �Z8��Q������j ������������PV�������6����������9��������*����?"u�� �������j|V�^  �����������������j"V�^  ����������t-1���������������эQ���������������I9��P���ǅ����   �A����E�x�t�������������������E;P�����������;P,�����������;P4�����1����������������D� �������U���������P�u�u�   ��U��WVS��  �]S������V�E�p�p�  S������S�U�r�2��  �� VSh�\������P��9��1ۋU��;Z}E�������QV�U�B�t��4��8
  ��Vh�\W��9��XZW������P��  C�U��;Z|U�B����  ����  ����  1ۋE;X4}E�������PV�U�B8�t��4���	  ��Vh�\W�Q9��YXW������P�  C�U��;Z4|E1ۋP,9�}���E�H0���8 u&C9�|�Q������Rh�O�u�P5���e�[^1�_�É���j"P�a\  1�1�������   �U�J0���8 ��t"�����<"��   ��5����G��F�< u�������Ƅ.���� ��W�4��  XZj �U�B0�4���[  ����t5P�U�B0�4�h�\W�`8��^XW������P�  �E���P,�)����v P�U�B0�4�h�\�ɍv Ƅ5����\FƄ5����"�c����U���B0�4�������W�  �E���H0�V����E�p(�p$h]������W��7��XZW������R�  ���:������2���Q�E�ph	]�ǋE�@ ���$봍v U��WVS��(  �u�4������t5�5��j4jh@[�y7���5��j.jh�[�e7��������e�[^_�ËE�     �U�E�    �     �U�����P�u������h   V�5����������tA���#t�X7��� ��f�P%   f��u7��-t2��+t-V�uh   W��4��������u����u��3��������^��������1��������р|�
�[  ������S��h���Wh�\V��5����H�   �E�    �<|t ��t�F�<|t��u����u�V3���������t�~ t�F�<|t!��tF�<|t��u����u�&3��1�������t�~ t��j|FV�qY  ����t(�U��<|t��t�F�<|t��u�뵄�t��~ u�멊��t��Ѓ�%�9  ��%�  ��#tZ��V�1  ����~�U����5������f�A%    f��u���P���F����E����~ �;���F���u��/���QWh]V�4��XZh]W�J  ����uP������Ph�sW�l4����Htk��h]W�  ����u2�E� �����S5������f�A%    f���l����������F��S������PhvW�4����Hu��U�   볋E�     먃�@��������n����~ �d���F������U���4������f�A%    f����������3���F�ސSWh�\�5���0��[�������������D� ������U��VS�]����u�  �C����   �C����   �C����   �S��u7�C��t$��h��P�B  ��h��h]V�0����1��e�[^�Ív �C��uɅ�t��jl�GG�������C��   ���sP�  ����x���s�s��  ���s뚃�h]��L��������RPh7]V�/�����M����v QPhB]V�{/�����*����v RPhK]V�c/���������v QPhT]V�K/�����������h�[�FL����U��WVS��(  �u��/������t5�5��j4jh \��2���5��j.jh�[�2��������e�[^_�ËE�     �@    �@    �@    �@    �@    V�u������h   R�������M0�������������   ���������#t�2��� ��f�P%   f����  ��-��  ��+��  1���������������ы������D
��x�
��  �������]]�   ���v  �������c]�   ���=  �������i]�   ���  �������o]�   ����   �������w]�   ��t;S�uh   ������R�M/������������� ������u�A.��������������������������  �U�B�$l   �D���U�����B��   ���U�rP��  �����s�����聚  �$�YJ���E�@    �@    ���J������������������  �U�B�ۍv ����������������
  �U�B뻍v ����������������
  �U�B뛍v ���������������
  �U��y�����@� �H������u�(-��1��u�����h@\�dI��U��VSP�]S�u�v�6��  �C@�������ك���u>�C8������Eu*�F�C(������u�C0��������Eu�   �e�[^�Ð1�����������U��SP�u�u�]h}]S�/���$�W  1��]���U��WVS���}�?"��t1��j W��R  ������t��)��e�[^_��1���������эA���B�B��u���j"�GP�R  ���x�\��tU���v ��j\R�qR  ������t�9�w��B�r����t<"t<\t���Ѐ: t�v ��9 ��t�B�J��v K�ݐ��j"CS� R  ���x�\��t�뒍v U��SQ�]��.�������f�A%    f��u��tC��1�Z[�Ä�t��C���E�t��.����E�f�B%    f��t�}� t	C�C�E��ߍC�����]U��ES��B1ۃ��Mt\��~G��t2��������Eu���ػ�����؋$�Ív ��������Eu�   ����؋�@$�B$��������u��؋�@�j��؋�@ �j �U��E� �P8�E� �@8� �*������1���Eu���ع�������Ív ��������Eu�   ���U��E� �@0� �E�E� �@0� �E��])���U����u�uh�6�ZN����U����u�uh�6�N����U���h�]h�6�u�u�q  �Ív U���h�]h�6�u�u�  �Ív U���jh�]h�6�u�u�  �ÐU���h�]h�6�u�u��  �Ív U����u�uh�6�vu����U����uh�6�u���Ív U����u�uh�6�Fu����U����uh�6��t���Ív U��WVS��<  �S���^_Ph�\�E����������   ƅ���� �v S�uh�  ��X���P��)��������   ��������W������S��H���Vh�]��X���P��*���� H��WSVh�]��X���P��*���� H~���������P�uS��  �����t�����������P�uV�/  �����T�����W�?  �<$�o  �U����   �e�[^_�ø�������P�p*����    ��� �����U��WVS��,  �Eݝ�����]�u����ZYPh�\�cD��������j�WVS�C  �� j���h���S�������������^  X�E��tPWSh�]�u��&���e�[^1�_�ø�6�ߐU��WVS��(  h   �u�>���������ܮ��P�Í�����P�v�v��  �� S������S�v�6��  �}�����H  ��������PWSh�d������1���)���� ;^}P��Q������P�F�t��4��E���������PWh�d������P��)����������P������C��  ��;^|��}����  �F����  ��xJ��E�]���F ���$��6t��]PWh�]������P�Z)����������P�������  ��1�;^4}e�v Q������P�F8�t��4������U�������҉$��6t��]PWh�d������P��(����������P������C�*  ��;^4|�1ۋV,9�}��F0���8 uC9�|��������e�[^_�É���P������P�   YX������P�F0�4��  XZj �F0�4���K  ����tN�M���F0���4���6t��]PWh�]������P�E(����������P�������|  ���V,�d�����U���F0���4���6t��]PWh�d밋U�����v��6t��]PWh�]�x����d�9����u]������U��WVS���u���1���������Q�T;����XZVS�M(���e��[^_�Ð��U��E�8 t�@�8 u���U��M�U�v ��AB��u��E�ÐU��UJ���S�M�]t��J�CA���u�� �E[�Ív U��UJ���S�M�]t���t�v J�CA���t���u�� �E[�Ív U��M����Ut��A�B��u��E�ÐU��UJ���S�M�]t��J�CA���u�E[�É�U��S���]�uS�����$�����؋]��É�U��S���u�]�uS������$�����؋]��Ív U��V�u��S�]ti�۸   tT���tD���t5���ЍA�FC��w�� �B���w�� 9Ѹ����|!#���t���u˄Ҹ   u
�; ����H[^�ø   �������U��WVS���}������1���ыu�y����t9�U�8�t�v F���t&8�u���tPWV�u��#������tF��uǊ   1�����H�e�!�[��^_�Ív U��WVS���u1������������Q�"��������t��VP��%�����e��[^_��U��SQ�E�M�E�����]��t�v 8�tB���u�Z��[�Ív �E����U��S�]��� �ى�tN��	tI9�t��@A��t���; ��t�@�8 u�9�tH��� t��	t	�@ 1�[��H��� t���	t���@��� t���	t�먐U��WVS��$jj�!���E�XZjj� !��_�5���E��!��^�5���� ��� ��������ts��xO�]�߉���S�}���$����9���t.@u��E��������u�j� ��XZ�u�j� ���E�e�[^_��@u����5��j&jh ^��#�����E�����뷃�j j�X ��Y[j j�M ���$    �uh QhQhQ�����j�5#���U����I���$�   �Ív U��WVS��  �u��~p����X���P�j   ���������������v ��PVh�^W@���0#���^��PW��X���PS�5  ��j S�Q ������t�S�9����e�[^_��������U��V�uS�.tmp�F �V  ����t�8 u��V�u^���e�[1�^�Ã�h�^V�N!��XZSV�E!������U��E�@h    �ÐU��S���]�uS�Ջ  �Ch   �]��ÐU��S���]�uS赋  XZ�u�C4P觋  �Ch   �]��Ív U��VS��  �u������QVh   S� ������tAP������Ph�`S�U!����HuӀ�����#tʃ�S�u�  ��������H�e�[^�ø������U��S��  ������S�u�'   ���������xPSh�O�u����1҉Ћ]��Ív U��VS��   �u�]� �Ch��~����x���PS�=�  ���������u�Ch��I��t1��t�   �e�[��^�Í�����P��x���Ph�_V� !�����ԃ���x���PV�!���鐃�������P�C4P�͊  ���������u��Ch�U��WVS��  �u�]V�,�������ɉ���   �ȍv </tDB���u���S��h���S��  ���������t
�e�[^��_�Ã�SV��������   ��v ��t�������9Ӊ�tC�@9�t�����  W������W豐  C����t�����롃�S��h���S蒐  ����u�PSWV����듊�U��V�uS�]�    �Ch��~��S�u�@�  �   ���ChH	�e�[1�^�Ã��C4P�u��  �   ���݉�U��WVS���u�u�}�Uh��������tX���uP�����É4$�n�����۸   u
�e�[^_�É��OZ��PW�u��h�^h�:��X����P��8����������#Z��PW�u��h�^h�:�X����P�8��������U��WVS���}W�]S�uV�@����1҅�u�e�[^��_�Ív PWSV��g��������tK���uP�����É4$������ۺ   t�W�u�u��h _h�:�/X����P�8��������W�u�u��h`_h�:�X����P��7��������j����v U��VS�Ā�uVh�_��x���h�@S�2��XZ�uh�_S�uVh�_�	����e�[^�É�U��S��   �uh�_��x���h�@S����YXh�_S� ����]��Ív U��VS�Ā�uVh�_��x���h�@S���XZ�uh�_S�uVh�_�����e�[^�É�U��S��   �uh�_��x���h�@S�q��YXh�_S�����]��Ív U��VS�Ā�uVh�_��x���h�@S�:��XZ�uh�_S�uVh�_�����e�[^�É�U��S��   �uh�_��x���h�@S����YXh�_S�(����]��Ív U��VS�Ā�uVh�_��x���h�@S���X�uh�_SVh�_������e�[^�É�U��VS�Ā�uVh�_��x���h�@S�~��X�uh�_SVh�_�����e�[^�É�U��VS�Ā�uVh�_��x���h�@S�>��X�uh�_SVh�_�u����e�[^�Ð�U��U�<.tB��t'�<.u��ъA���Rt�<0t�J�ȉ ��u�� 1��ÍB�쐐�U����,���t�Ív ������$�������t-���0��������,���u΃�h�O������,���뷡,��ސU����}�E�U�Mt��QRP�   ��1��Ð��QRP�]F  ��v U����}�E�U�Mt��QRP�P   ��1��Ð��QRP�uF  ��v U����}�E�U�Mt��QRP�   ��1��Ð��QRP�F  ��v U��SP�u�u�]h}]S����$����1��]���U��VS�}�]�ut�u�]�e�[^��  ����VS�JI  �����   t	�e�[��^�Ã�VS�w  ��1҅�t����`����1���u��`��������u��   ���뵍v U��VS�}�]�ut�u�]�e�[^��  ����VS��H  �����   t	�e�[��^�Ã�VS��   ��1҅�t����;��������E��uj��� 8�����������E��u���������������`������Eu/� 8������������E��u��������������   �k�������������붐U��WVS���}�}�]t3��SW�A   1�����t�����������Eu�   ��e�[^��_�Ã�SW��G  �����   u��U��SP�E�U��E� �     �@    RPh�`�]S�����Ht
1҉Ћ]��Ð�}� u��; t�C�; u��K��A�1�<vڍA�1�<���ΐ�U��WVS���u�  ���������������x��t�e�[^1�_�ÐJ�E��s  �E荘t��t�����P��+���=x��������  �������  ���������������(7����ܠ,�����1ۋt�݀�������9������^  �}�x�f�E�f�E��m��U��m��E�������Eu�M�E��x�E�;��   |�E������E�@�C�t���9���|��؋=x���tP�����ى��������� �����D��������\�����������l�����\�����ˉ���������% 8ܠ,�����1�����9ˋ���ܰ�}i�}�x�f�E�f�E��m��U��m��E�������Eu�M�E��x�E�;��   |�E��������u�E�@��t�C��9���|�������������������������E� �� 8�D������������E��ud��������D��v ����������Eu�������ډ��������,�������Eu�������������Et������������������������Ã���t����  ������x����U��E�@(�e�p �Ív U���E� 8���E������������E��uA������������Eu����v ������������u�������������t������������������Ӎv U��S���]�{�Et�]����sD�s@���$�k����C8�������ك���Eu��C@��� 8�������ڀ�E��@u�����봐U��S���]S�u�u�����c@�s�]��Ív U��E�@ �M�h(�Ív U��E�@�M�@@�Ív U����   �p��É�U����	   �t��É�U��������t1��Ð��hh����   �B������U��WVS���E��E�]��������M�DQ�$�D�}�f�E�f�E��m��U��m�]�$�$��������E�   uKA�5p�9�}V�E��E�U����݀ �݀���v Q���$���m��U��m�U�$�$��������EuJ9�uAG9�|����؃�[^��_�������𐐐U��WVS��  �]��~P��   �   w��N�����������t
N�  @���u���~%����   �   w��PVW�u)���������ݍe�[^1�_�Ð��U��WVS��   �5���}�]��x����a���������5��W������5��jjh@a�������x ���۸Gat�LaP�5�����������5������4$�*  ����t���V�I�����x�������Yt��Y~��nt��yu��   �e�[^_��1����u���d��������Nt��V���U����uj �u�}����1��Ð�U��VS���M�ɋU�]�'  �B ���������	  ����  �B����������  �r���3  �B(�B0������u,���؃�t�E�a�E�:��[^���J���E�a���B8�B@��������   ��u>�B �������}������(7f�E����f�E����m��]��m��E����Bu�B   ��u>�B�������}������(7f�E����f�E����m��]��m��E����Bu�B   �J��x<�B��x!��P�����4$�Z ��$�4$�Z��[1�^�����������E�a�
����������������������E�a������B(��`����������Etf�B0��`������EtD�B8�B@������u,� 8�v �������������R8u�������������p��������g��������E�a�p������E
b�b������E%b�T����B�������EBb�=�����ETb�0����r��������Eqb�����U��E��tH������   ��P���1���U���jP�����@�$�1#���Ív U����u����YZPR�����@�$�#���É�U���jQ����@�$��"���Ív U���jP����@�$��"���Ív U���jP�v���@�$�"���Ív U���jP�Z���@�$�"���Ív U���j�u�   @�$�"���ÐU��U�Ҹ����~������t@��U���j�5h�j �u�u�u�u�  �ÐU���j�u�u�u�u�u�u�]  �Ív U���j �5h�j �u�u�u�u�7  �ÐU���j �u�u�u�u�u�u�  �Ív U���1��} ����P�5h�j �u�u�u�u��   �É�U��1��} ���M�U ���E �U�M��   U���j�5h�j �u�u�u�u�   �ÐU���j�u�u�u�u�u�u�y   �Ív U����`���u���u�r����`��d� 1��É���P������Չ�U���h�ch�:�F��ZYPh �����`�����u� ��Ív U��WVS���  �u�=�����5���^	�����=d� �8  �`��ɋU�d���t�E��t�E�8 u�E    �E�  �E��t�E�8 u�E�E��t�> uC�} ��  �} ��  �} ��  P�uh�ch�:��E��^_P������V������G���������������SVh�c�5���F�����uh�bh�:�}E��ZYP�5���#���]����th��h�ch�:�SE��ZYP�5�������E����t�E�8 ��  ��hdh�:�E��ZYP�5������[X�5��j
�	�������A�����Phdh�:��D��ZYP�5������5��jjh=P�4����W�G#  ����������W������Wh%d�5���C���������� �1  P������1��} S��PW�  ����v�5��jjh+d�
���������$��d�5h��] �ۋ����u��6P�u�u�1  ��Q������S������PW��I�������������  ��������P�C�����������U  �E ��ukPh�6W�u�S+��������u$QWhBdh�:�C��[ZP�5���G���C����������t��������P�u�
�����؍e�[^_�Ã�W�勅�����t-��S���������������   ��������PW�?
����P�����W�u�*�����} u���U�����W�u�
�������놃} ~K�} ��   ��t؃} u�PWh ch�:��B��Y[P�����S�	��XZj S�/�������� ���뛃} ��   ��t�PWh`c�����PWhYd�����RWhvd�������W�����u�)����5h�S�0����u��1�������v SPh�d����P�uh�c�W����E ���>���P�uh�d�?������5`������`�    ��������h�dh�:��A����P�!���v U��WVS��   ��h���P�E�P�E�P�u�Vh�d�u�E� �E� �E� �P���� 1Ʌ���~=�   �d������1�8�u$���   t��������}�-t*�������t
�e�[^��_�Ã��E�P�u�O���   ���u�������tԀ}�ft������ǀ}� u���   t����E�P�u����   롐U���X��������}���É����$B��ZYPh#e�3  ��������1҅����~�P�E�P����A��ZYPh#e��  ����x"�?V  9E�t���    1���_���9E�u���5����  �A��ZYPh#e��P���������x���   �   �L�����h eh�:���    �@����P� ��닍v U��������~���5���  ����������������1���U����=���|1��Ð������������ꐐ�U��S���]�C    �C
   h�   �����C    �   �]��Ív U��WVS���M�ɸ   ��   �U�R�E� �҉E�U���   �M����E��M���M�Q��H������t�U�E�@����E��U�M�ԋU��~R�U����E�   ��  ��������)��5���U��������u�E�V��P�s  �E��@    ���M�E�M��~2��U���M����Q�E��U�6H������t+�E�@�E�M��ϋE�U�M�P�1��e�[^_�Ív �U�����   ��������)U�   ������]�Ë9�����   9���   �S��ۋU�E�B9E�}EP�E��u���E�VP�E��   ��93~�ߋM��E�y�C�W����C�U��M�B�K�C�����
���B��P�u��+���E�����]�Ã�딐�S�y����C�M����������g����������։���)�J�#����������։���)�J�k�����U��VS��j�t�SK�u�n��������Ft�v K�     �����u�E��V�E��   �F    �e�[1�^�Ív U��WVS���}�E�    P�u�~F������t�F��������e�[^_�É��^��~5�U��xD��������)U�   ������9�t9�~�D���1�붋D��D�U���뚉������Ӊ���)�J뵍v U��M�A��~,�A   ��B��t�v �A���D��u��A����1��ø   ��U��S�]�C����D1Ʌ��Ct#��x&���D��t��C���D��u�   �ȋ$���؉C��v U��WVS���]�C���}~j���KA;t��K}>�S���3�D�����t܋��x��ȋU��   �e�[^��_�����D���S�B�����1҅�t��C�����1���U��E�P�E�ɸ   Ív U��WVS���}�   ;w �   �����tF� ������;w~���7� ���e�[^1�_�Ð�U����U���   w/����Ѝ�������~Ht��jR�  �É��U��R���������U����U���   w/����Ѝ�������~Ht��j R�`  �É��U��
���������U��WVS���E��E�U��1ۍ4 �p������3����  C���������~�E��E�U���<�    ����p���   �������   ������   ����t����  �r���X���  �f���^���  �Z�����l�Y���  �H������  ����u\���  ��Ǉ������u���u������e�[^�   _�Ã���x�P�<�����<��P����tɃ���8�P�҃�븃���4�P������됃����  �������/����U��WVS��C  �E���{  �E��E�U����    ��h����   t��t����   9��  ��  �E���UE��V������l����  h�H��d�����x���P������9��Ph�Y��x���R������P�  ����x���R�K:���������$�=������  �����H  ���u��A  ��`�����`������ɸ������  ��t�;��  }H��d����≕\�������u������+�t�S�\����4�P���`���C�B  �� ;��  |ǋE��E�U���4�    ����t��t���l����   9��  �  ����`��������XZ������P�E��E�U���4�t����  �*��������y  �����  �!������E��E�U���4�    �����  ��p���l����  ���i  ���u�  �����+  ��h�H�8��XZh�  P���  ���  h�H������P��  ��P������$�����`�fcelf�d�l �����u������E��E�U���4�    ��h���t����   ǀ�   �������  ������h����m  ���  ���D  �E��ǅl���   t��p����  ���u  �E��E�U���<�    �� ����@  �M����   �]���E]���4�    ����,��H���X��0��<���1�����p��������  F��������~�E��E�U������    ��p�������������u��l����e�[^_�Ã���x�P�������ރ���l����  �H  ��������Sh�_���  �  XZS���  �  ���  �����  ������P���  �̙��[���  �`����E��E�U������l����  ������  ǂ�   �����E��E�U����    1���h�������p������   ����P��l����  ��-  ���  �����  ����x�S謅����S���  ���  �ߒ��������   V��t���S��p���P�E��E�U���<�    ����P�����$�O=������t
ǅt���    S�����Sj ��t����	Z  ZYS��l����  ��U  �$�M[  ���  ����u
������u&�E��E�U�����4�,���  ���t���������S���  ��  �$������ك�hHf����������P���  h�H��x���S�4������  hafS������S�  ��S�����뽋��H���   �>���������P���  莘�������$�|����������P�.������������  ��,�h`�������V�
  �4$�Q���[XV���  �3�������x�����  �.������;���V���  hif��x���S�^����$������������V���  h`e������S�3����$���ǅl�������롍v ��P�s���ǃ�      ��������P�X���������Q���  h�e������S������$�d�����������  ���  h�H������R�	  �������$�M��������  h�H��x���R�������  hI��x���P������R�Q	  ��������P����X�u�`�cell�d� �l����r�����p����  Pjj R� ���������X�u�J  �������������P���  hif��x���S������$���������g���������R���  h�e������S�����$�C���9�������x����   ��p���X�����<�����  ��;��   �������T�����X������u���   S��T�����p���`���C�X:  �� ;��   |��r�������$�������������$��������l����  ���  �E  ���  ��;��   }"�P���  ���  �uC�R,  ��;��   |ߋ]��]�E������t����  ����ǃ�      �������U��WVS��  �u���������l����  ��u��h f����1��e�[^_�Ív �;*�����  ����   PWh1Ih'Z�S*����Whrfh>I�@*����������4�    ������t]P��,�h�H��x���S�������0�hIS��x���V�  ��S�r0������t���PWV�,���<$�M,����t����C���P����h�s��x���S������WShvf�)�����t����v PWh8I�+���U��S�]��K���M�U~����BAK���1�[�Ð�U��WVS���   �����t�   �e�[^_�Ã�hzz���   ���    �D  �����Ǎ����tu�PWh�   V��#������tT���������tD<:t	C���u��ӄ�tσ�V� C�����$�������> t��; t���SV�   ��랉���Ń�W�c�����1��L����U��WVS���E��t�8 u���u�  1��e�[^_�É���P�k����$�E��(����E���8 ��   1����9��E�����}�=��������   �u�F9�|�u���x(���u��������U��ӋM졄��L��v����C�ۉޣ��t:����P�5������Y����u����������U졄��T��.�����j����̉����uP�|��������_����E�D��   �������P����_�u�   ��U��WVS��1��=��9�}-����E��v �E�����t���uS��������tF9�|�1��e�[^_�Ã�S�7��������    �   ��U��WVS��1ۋ5��9�}&�=����߅�t���uP��������tC9�|�1��e�[^_�ËD���U��WVS��jj�����[^jj�E���������$�q�   ������t31ۡ��9�}������څ�t�L���u3C9�|��V���������u�j����XZWj�����e�[^1�_�ÐQ�E�Ph�`�t��)�����Ht���뭡���t��4�hE;V��������U��������t���uP�U����Ív ��h�f������������uփ�h�fh�:�*����P�	��U��S��@�]S�4   ����t�]���PSh�fh�:��)��ZYP�]�S�#����$�{	���v U��WVS���]�޿�>�   ��u��[^_��_����v �����]��[^_�����U����������u�u�W����B���1��É�U����q������u�u�3���1��Ív U����Q������u�R�������1��ÐU��������u1��Ð��������U��VS�]������x*1ҋ��9�}�5����օ�t�8 tK���tB9�|�1�[^�Ív U�����    1��Ív U����E�����    t�8 u1��Ã�P�����������U�塘��É�U��SS���������1ۉЉ��1�9����    ���    }#�v ����Ѕ�uC;��}�����v 1��]��Ð���t��4���������С��U�������壄�������������1��ÐU��WVS��  �]�u�(���ǋE��t�E�8 ��   ��t	�> ��   ��(��PWh�@S���������W�)���E����t�E�8 u;�M��t�E�8 u�e��[^_�É���h�^S�"���XZ�uS�������։���h�^S����^_�uS�������막�V�u�����P������P������P�u��,�������>�����������P�u�����������PWh�@S������ �3����U����u�uh�H�����U����u�uh�H�Z����U��VS���]����؍��4�����xL����؍�����p����   ��u�؍e�[^�É�������j@P�N �����  �$�H   �Չ�Qj�E�PS��������t����؍�����    눀}��u�}��u݀}��u��q����U��WVS���u���������    ��p��E苀�   ����   Pj�E�PV�G�����HtE�������W����0���,���h�gh�:�A%����P�0��������e�[^��_�Ð�E��t���t��]䋛�   C���؃�S������SPV�E���������9��z����U�1ɋ��   9�/�E��u��1��E�9�}������GKu􋆀  ��A;M�~ك��u��b����   �a���������   PS�U����  V�J�����9غ   �3���������U��WVS��j j �u�����E��E�U���<�    ��t����   ��   �$�E��'����E�� �M�1�A��;��   6��p��}�ߐ�U苂�  ���   �؈��K���F��;��   ~�Q�u��u��u����Z�u�1�;E����n����e��[^_��U��WVS��  ��h���P�E�P�uV�}W�(���������������d�����  P��h���P�E�Ph�Y�2����������   Qj�uS蘑����`����$�z�����`�����1�����   VWh�gh�:�#��[^P��h���S�W�����1���������эt���d�������td��h���W�E�Ph hh�:�"��_ZPV����ZY�1��߹���������`����t�V����X��`����I����$�u��������e�[^_�Ã�h�h�VWh�gh�:�U"��Y[P��h���S�������1������򮍅h���P�}�Wh`h��h�:�t��"��_ZPV�u�����1�����������h���P�}���W�t��X�������u)��h�hh�:��!��ZYPV�.�����h����$�:�����h�h�Չ�PVWh�Y�1���������V���VWh�hh�:�!��[^P��h���S�����������U��WVS��   j ���    �'���������`���u~P�5��jd��h���S��������ƹ����1����Ƅf��� Y_S�u�"�����`�������u!���   t�e�[^_�á����tR1���v ����d���j��������ʍv ��h,�j����������d����b�����Pj�������O�����j�����v U��S���]j S���   �`���XZSj ����Y[h��j�H�����XZjQ�l����$����XZSj�*����]��ÐU���Ð��U���h`i� ����Ð�U��E�     �@    �1�ÐU��WVS���   �}W��������uh�H�����V�4������uhfjV�W������u0�u�uh�ih�:���ZYPV������4$����1��e�[^_��P�uhfjV��.����������   PSh�   V���������t{�����P�����PhpjV���������uPW�����������  ��볃�W�"  �$�b����u�uh�ih�:����ZYPV�T�����V�����������M�����S�(��������u!�u�uh�ih�:���_ZPV����[뽃�W��  �   �����u�uh j�ʉ�U��WVS���u��  �ǃ��������t,�E1ۋ9Ӌp}�v �D���uC9�|��W�����   �e�[^_�ÐP�4�hxjW������E����ˍv U��WVS���u�s  �ǃ��������tP���u�����u����]�P�uVS�%�������t�E���~�P�u�hxjW�p������Ӄ�W�����   �e�[^_�ÐU��WVS���]S�z���X�u�A����}����u�P�uWV��������tPS�u��u��a  ���܃�S�   �e�[^1�_�ÐU��E� �É�U��U�ҋEx;|1��Ív �@����U��U�ҋEx;|1��Ív �@�D���v U��SP�]���~���s�������    �C    �   �]��ÐU��WVS���E����   ~(�   �U9ًz}�W���9B�}A��9�|�   �e�[^_��9�}�h��jSW�   �����1Ƀ�9�}!����9�E�t!���D��BA�E��F9�|�A�U�1�뫋D�B���U��E��E� 9¹����|1�9������Ív U����M����   ~h�jR�q�k���1��Ív U��VS�u�]�K�V9Ѹ����|9Ѹ   ��9Ѹ����|1�9����[^��U��WVS�Ā�}Wh�H��x���V�����[XhfjV�*��������t
�e��[^_�����PWh@jh�:�@��ZYPV�����4$�'������ʉ�U��S��x�u�]�h�HS�t���XZhfjS觝��1��]���U��WVS���]1��9ȋu�}}�S�v 94�t@9�|�QSWV�]   1��e�[^_��|��   ��U��WVS���]1��9ȋu�}}�S�v 94�t@9�|�PSWV�   1��e�[^_�É|��   ��U��S���]�@���P�s�������U�T����U�C�T���]�1��ÐU��U1��
9�}�R�v �D�    @9�|�1��Ð��U��WVS��h$  �}W�Y������u�uh	k�F)��������t!QPjPW�#������u@��t��S������P�u�u��h�jh�:�����P����������e�[^_�Ð��W�G/  ��SjP�wPV��������t���V�(/  ��SjP���   V��������{�����V�/  ��SjP���   V�|�������U�����V��.  ��SjP��@  V�V�������/�����V�.  ��SjP���  V�0�������	�����V�.  ��SjP���  V�
�������������V�j.  ��SjP��0  V���������������V�D.  Ǉ�      ���  ����1BR��S��jP��8�  P�������t$���  ��������8�  P��-  ���  밃�S�m���1�������U��WVS���]Sh	k�'����������   P�uh�OW�����E����PPh�OW�|����E���   Ph�OW�e����E���   Ph�OW�N����E��@  Ph�OW�7����E���  Ph�OW� ����E���  Ph�OW�	����E��0  Ph�OW�����1��E��;��  })�ÁÄ  ��PSh�OW�����F�E����P;��  |��W�P���1��e�[^_�Ã�S��h�jh�:������P������������U��S���]�-A  ZYPS�����YX�u�CPP��������YZP���   P��������YZP���   P����XZ�u��@  P�����a����Phkh�:�U��ZYP��0  P����ƃ�   ƃ�   ǃ�      �   �]���U��MS��ҊEt8�tA���t8�u�����t1������X�!ˉ�[�É�U��US�1ۄ��Mt��8�tB���u��ɉ�t��[�É�����U��WVS���E��E�U��j �4�8�V�F�P�]K������E�    �E�    �}�t�v ��WV�>�������tKK���u�1�;]|�   �e�[^_�ÐP�uS�u�/  ��@tC;]|��׃�Sh@k����������ǃ�Sh�k��U��WVS���E��E�U��j �4�8�V�F�P�]K������E�    �}�t����WV�F�������tHK���u�1�;]|�   �e�[^_�ÐR�uS�u�  ��@tC;]|��׃�Sh�k�o���1��ʃ�Sh l��U��WVS���u1��1�9�}���F���8 uC9�|��e�[^��_�É�P�F�4�hE;�u�������@����H	ǋ�ʍv U��WVS��  �O����1���tl�������P�uh   V�1
������tj����������tZ<:tP��C���tA<:u���V� C�����$������WSV�%������u���W���1��e�[^_�Ív <:u�뽰:�����������U��WVS���u�V�}W�*���ËE�����t
�e�[^_�É�RS�u�u�������u��S�'���������PVSW�{���$����E�뼉�U��WVS���]�E��}� P�u����ƋE�����t
�e�[^_�É���V�u�t������t)QWPS��������D� �E�   ��V����E�뽍v �E�    �搐�U��E�ԏ1��ÐU��WVS��h�j�u�Ļ    �F����}�����E��E�    t�E�8 u�E�E��j����������M  �=��Wj/jh�l�z�������t	�> �
  1ۋ5Ļ��uT��S���������t���uV�u�uW�=  E��� C�ȡĻ��u�]�����   Wj/jh�l������;=��t��W�u[�������u�j�i����ԏ����u
�e�[^1�_�Ã�j�(�������t��hmh�:�;��ZYP�5��������������5�����������
u��Q�uhmh�:����^ZPW�������D������uV�u�uW�Q   �E��� ������h�qh4m��Y�������������������U���h��u�Ļ   �����ÐU��WVS��<  �}1��?.u
� ��  Wh�6�u������S����XZj S����������v  �E����  PShAm��h���P����Y[hzz��h���P�!Y���������8  �Ļ���  PSh�  ��h���P�D��������  F��t{�E��u���u��h���P�*�����뱀�h��� ��h���t��h���<
t=B���u�P������PW��h���P�U������P��h���PhHm�u������ �[���� 뾉�W�uh�lh�:�A��YZP�u������U�����`���P������PW������Pƅ���� ƅ���� �U�������� �(���������P������PhGm�u������������S�X�����Ļ��u��~���uj
�b������e�[��^_��PShVm�i����������!����U��E��� P�E�P�E�P�E�P�u�u�  ���E�P�u��u��u��u��u�   1��Ív U�帀m�É�U��E��� P�E�P�E�P�E�P�u�u��  ���E�P�u��u��u��u��u�c   1��Ív U�帎m�É�U��E��� P�E�P�E�P�E�P�u�u�g  ��j �u��u��u��u��u�E� �   1��É�U�帝m�É�U��WVS��\�u�uhv�u��EV�}�]�E���������E�Ph�OV�����E���m�������ك���u��C��;�E�    �E�    ~1�G����m������E��   ���$h�mV�i����4$�A����E���<0u�}�0u	�}� t3�v <0u�}� t&���E�PVSWh�m�u�&����� �e�[^1�_�Ð��~���E�PSWh�m�Սv ��~�E�PWh�m�u�����������h�m������u��u�hv�W�����U����E��������E�Uu!���S���u�u�u���$�   1��Ð�N�ߍv U����E��;��������E�U��   � 8�����������Eu����v ������`������EuQ� 8�v ����������Eu����v ������������Eu ���W���u�u�u���$�   1����E���������U��VS���E����������E��@�M�u�]u���    �    ���[1�^�Ív �}�f�E��f�E��m��U��m��E����P�$$��m�����m��]��m��ɋU�����H!Љ�!�ɉ$�$$���������Ƀ���E�t���돐��U���jZ�uh n�u�T   �É�U���h�   �uhn�u�5   �Ív U��S��x�uhn�]�S�����j �uhnS�   �]��Ív U��WVS��,  j�uh�m������P��������x���Q��X���P������W������S������Vh
n������Q������ ����  ����x���PWSVh&n������Q������ ���x  ����x���PSVh)n������Q�l����� ���F  ��x���PVh,n������Q�G�������t1ې�e��[^_������ǅ����    ǅ����    ������1ۅ���  ������1ۃ�;��  ������1ۃ�;��  �]����  1�;E��  ;E�P  �م��  ��t.��������Pݝ�����2  1ۃ���݅������   ������Q��m���$��ڽ����څ�������5@n�����M��x����P�����M�����������E����@u��x���<�   tg<@~<Z	�� ��x����M�8�t:At	�����������y���t	��������8�t���ػ   ���������ـ�E��@t	���M�����������������x�������s�����������Qݝ������   1ۃ���݅����t��������������=�����~	�����-�����~	����� �����������E��������
���������������q�������������v ��������������������������������������X���������8n��X���t)��m����0PB����$��������u�����������������U��U�<:tB��t/�<:u�B���01�<	wB���01�<	w�B��01�<	�����ù   ���U��U�<:tB��tC�<:u�B�<:t��B��t/�<:u�B���01�<	wB���01�<	w�B��01�<	�����ù   ���U���h�   h��� �����_� ���Ð�U��VS��  �uVh�Y�;��������tPj�uS�  �$�V���1��e�[^�ÐSVh�nh�:����ZYP������S�<����$�����������ɐU��E��x�����������É�U��WVS��T  j �}W���q��  �����������   ��������4�    ��l����  ����    ��   ����x����   �5��蒹��XZ�5����   j ����uW�o  �� ��������ti���   t`���������    ��h����  ��������uC��x�j����P���   �u�l�����������  XZ�5��W�  �e�[^��_��Q����P��x����   �u����������  �5�h�n������S�����$�����U��VS��j�uV�]���q�  ���������u�e�[��^�Ív Q�EP�EPV�  ��XZ�5��u�u�uSV�F  �� ��������t����   t���������4�    ������uP����P�uS�Xk���   �P����P�uS� ������ҍv U��S���]����؍��4���uS���q�  ����������t���   t����؍�����   �Ћ]��Ív U��WVS���E�]�E��u���qj S�Y  ���������th����؍��<�    ���9��5���   ������    t_Nt@��t5H������   �u�S�� �1҃��=� �T��e�[^��_�ø   �҅�tH������   뾸   뷐��tH������   �1�랃���x��E����   �5��臶����Vj �E����   j ����u�S�  �� �����   ���   �e�������   ����؍��4�    ������uG��x�P����P���   �u��_i������؍��������E�]���e�[^_������P����P��x����   �u��������랉���؍���V����R�����u��i��돺��������U���j �u�u������Ív U���j�u�u������Ív U���j�u�u������Ív U��WVSP�E�E��E ���}�u�]�MuX[^_��!��E�E��M�]�u�}�EX[^_���  �U��WVS��,�E��E�U����    ��h����   1������E�u1��������}�E�x�E;���|
1��e�[^_�ËU1���~�u���Y  �E���-  �u�����tC�M���E�   �  �E��E�M������E��E�    �E9E���   �U�J�Uȉ����M��Q�E��o	����������  �U�1����E�    u�UUԡ����E����R  �E�    �M�1��ɋU�~�E�������tF�E����J���M��UЅ�t���   ;u�~�u��EԋE]�9E��^����E����  �E��E�U������h��M�;��  ~���  �U������}��U�wK����E�    �U�H9Uԉ�}7�   ;U�~JC;U����J��~������CAJ����EԋE9E�|Ρ���=���U܈�M܈��1��ECG9Ɖ]��E�    �E�   �E�    }^���   tP�u�S�u��  ����u3�U؋M܍T�E�9U���   ��PQ�u�GW����1�}܉]̃��EԋMF]�9M�|��E��t&��t�E؋U܍D�M�9ȉE�|b�E�    �E��uE�U��UBVR�U��5���u������;E�t���u�u��  ������P����   �F���W�E��u��5��뿉��P�u��u�GW�q�������E�    �\����E���ME���US���R�5���U�Q�t������E�   �E������E��������u���|����E����a����E�   ����Pjj �u�����%����U���������E����E���  Rj P�u��������������������v U��S��t�U����Ѝ����������Mc��|:�ɺ   u	�Ћ]��É���,��5�h o�]�S�����$�:���1��щ�JtP�5�h@o����,��5�h�o�Ń�uڅɺ   u���,��5�h�o뤍v U��WVS�E��u��1��ҋ]x%����؍�����9�~��)щ[^��_�Ív �����     1��͉�U��SS�U����Ѝ�����t����  ��t1��]���R�u��,���h ph�:�\�����P�K���ǃ�     �ȍv U��MW��VI��S�u�]~����CF1�8�u��I���   [^��_�ÐU��V�u�������S���P�]S�5��V�5�����9�t���uV�*���������e�[^�É�1���U��S���]����؍�����EP�5��S�T&  ����x	1��]��É����uS������������U��VS�]����؍��������u��U���Pj RS�{�������x1��e�[^�Ív ��VS�v����������v U��S��j�]j S�@�������ڍ������U���]���U��U����Ѝ����������Ív U��WVS���E��E�U����    ����1������E�1������E؋E���ux�E;���|1ҍe�[^��_�ËE1҅�~�}܅���  �M؅���  �E��E�U��������j ���R��8��5��W�ս��XZ�Gj W1��P��;]}�}�"  ��V�������t#�E܅��E�    �E�    u�Uڡ�����V���E��E�PW�U��{���������   ���u�i���ZYPVC�?c����;]��|��E��E�U����    ��<��H��u`�E؅�t9P�u�u�u������@�������������u�u�G������   ����P�u�u�u�������@�����������փ���8�P�у��P�uSh@p�����������b�����V�������t@�E܅��E�    u�Uڡ������E�PW�������������P�uSh�p롋�E��Ճ��u�u�[���������S�u�u�u�������@���������������U��WVS���u������������E썇t���   �E�B;E��   ����   ��V��   �E��U����Ҹ������   �U��x���}�1ۉU��}���   ;��   }/��V�M����   P�E���4�P��u��  �� ��xpC��~��E���~���u����������������t�P���������    ��t�)M�����U�B�4�P��u�*���   �e�[^_�ø�������U��S���E�����j ��t����  蔹������t�����  h�p�����������]��Ã�j���  �@����Ã��۸����~݁��   ���щ���h q�����$����볐U��WVS���u�}�u�9�����j ����PW褺������xQS�uW袷����9�t/��V��h�qh�:�1�����P� ���������e�[^_�Ív �   ��U��VS�u������������������J���M~���������J�������������E�u[^�����U��VS�u������������������J���M~���������J�������������E�u[^��X���U��� h@qh�:�C�����P�2�����   �É�U��� h�qh�:������P������   �É�U��VS���u������������������J���M~����������J������������4��V�����e�[^�É�U��VS�u������������������J���M~���������J�������������E�u[^��@���U���Ð��U��WVS��  �u�V�u�u�IS����1҅�~eW������W��x���SV�']���$�#�������u��W��������t;�u�uh rh�:�����ZYP������S� ����$����������e�[^��_��V�u�V�u�u�T����1҅�x�S��t���W��p���SV��[���$�#�������t��W��������u7P��t�����p�����������������|�����x����u��H���   �r����u�uh`r�<����U��WVS��
  �u�u��@��XZ�uV�z������u/�uVh�r������S�6����$�����������e�[^��_�Ív P������S������WV��������t���uS�������������u���W�uhis������P�ѷ��������PV������P� ��������t>���uP��   �ǉ$茶�������   �c����uVh s������P�w�����SVh�H������P�a������uhaf������P�J ���Ã��۸�Wt+���uS�X   �ǉ$���������   ������ss��P�uVh@sh�:����ZYP������S������S�v���1������v U��WVS��,  ������ǅ����    ǅ����    ��W�uh   S衴�������`  �޿ys�   ���@  �޿�s�   ���  ��������P������W������P������Vh�sS蒵���� ��u5P�������������������������������������u�AF���� �U�����u	P��������WVh�sS�:�������tSWVh�sS�%������������������������������������������u�=E��ǅ����   ���������������������������������������u�kD��ǅ����   �čv �E�@   �   �e�[^_�ËE�    ����u�C������~���u�F�������u�gC��1ۃ���~	�   ���V������V������W�u�FD�������QVW�u��D��������ʍv U��WVS��,�}����u��   �G��tVjjh�s襴���e�[^_�ÐS�E�P�E�PW��C������~���u��u��u�h�sV诰���� Q�E�P�E�PW�ID������~���u��u��u�h�sV������ ��W�B���Ã�Kx��v ���E�P�E�P�E�P�E�PSW�fB�����u��u��u��u��u�h�sV�1����E܃� 9E�tRPh�sV��������Vj
������Ky�����Vjjhys�����U��WVS��  ������S������P�uV�}��������t��WS良�����������ux�������>�����WP�h�������uiWVh�H������S�.���Y^hafS�ao���$�����XZhafS����������ú����t���uP�.����$�ڱ���   �e�[^��_�Ív PWhis������S�Ų��Y_VS��n���$�d���XZV띐��U��VS��H�]Sh t��n���}�����P�u�htV����XZSV�n���e�[1�^�ÐU��WVS��  �}�wVh@t�u蜮�����whPt�u������胮��VS�w,�w(誖����Sh`t�u�e���VS�w4�w0茖����Shpt�u�G���VS�w<�w8視����Sh�t�u�)���VS�wD�w@舖����Sh�t�u�������wh�t�u��������wh�t�u����VS�w�w�|�����Sh�t�u�ǭ��VS�w$�w �^�����Sh�t�u詭���U����u�e�[^�   _�É�P�7h�t�u耭�����wh�t�u�m�������U��SQ�]蟜��H���t�H�    �����u�Z1�[�Ív U��SS�v��������u�I�������J������Et
J�  @���u�1��]��Ð��U��E���dP��m���E���U��MS�����t�v �B�<^w�AC�����u�� 1�[�Ð��	u�� �㐐U����   �v U��VS��j�u�]S�uVh�u�  �� ���t9@t
1��e�[^�Ð��uPSV��h`uh�:������P����������Ή���W�ҐU��VS��j�u�]S�uVh�u�   �� ���t9@t
1��e�[^�Ð��uPSV��h�uh�:�:�����P�)���������Ή���W�ҐU��VS��$�u�V�u�u�1K�����������x(P�]�S�E�PV�bR���$��������t�E�    �U�e�[��^��U��WVS��L	  �]ǅ����    ǅ���������޿�u�   ������8�ǅ����    ��  P�u�uS������ƃ��������toPVh   ������W��������tqP������Sh�uW������H��  PShtjW�׭����H�i  �]��u"��V�]�������������H��!Ѝe�[^_��QVh   W�7�������u��V�'���������ԃ�W�'���XZ�uW�l  ����������x�U�B���������=  ǅ����    �PVh   W����������
  ��������tS�uW�������*  ���������Ív Q������Sh�`Wƅ���� ������HuՀ�����#t̋�������ƅ���� t%��S������P������Rh�uW詬���� ��tkS������PhvW莬������~��j �uS������RR�	  �� �^���S������Rh�uW�V��������������j�u������SP��R����j�uS������P���������V赫��1��b���PVh   ������S���������`���PVh   W���������H�����������P������P������P������Ph
vW讫���� ���������u�� م�����\$م�����\$م�����\$م�����$S�d  ��0����ǅ����   �����ǅ����    �x�������u�u�r���������������U����   �v U��E�@��u�`���U����E�E��u�E�P�   �É�U���j �u�u�5   �Ív U���j�u�u�   �Ív U���j�u�u�   �Ív U��WVS��t�]S�}W�u�7�������t ��hvh ��"���� ��e�[^_�Ð��SW� � �R��X�F �$P�]��}��4=���E��<$�5�������u�U�;}���   ����u�릋V�҉U�� �t��E��]��E����N�F�]��N�F�]��: � �t���<$��t�B�U�C�U��: u�� �O����B�U��A<$��   <?tIPW�u�V�E�P�  ����u�$���E����D���$V�u�V�+����E�����t���F�C��u���u��u��u�V�E��QP�U���  �E������l�����F�C��u��\����Q�$�M�����U��M1�;}���   ����    @;|�1���U���j �u�u�u�>   1��É�U���j�u�u�u�"   1��É�U���j�u�u�u�   1��É�U��WVS���]��K���u~g�E�x ���uV��P��X�$W�j;���M��$�E��h�������u/�U��E;9�M���   �����u�d���ZYPV�;M���ƃ���K����   �e�[^_�ø������v U��Eǀ�   �����1��U��WVS���u���   C�~ �E�    �E�    ��W��6����9�}*�u�uSV�c  �E����   ������uC���E�   �U�1���t���   ���E����   �E��e�[^_�É�U���j �u�u�u�u�   �ÐU���j�u�u�u�u�   �ÐU��VS���u�E�P�E�P�u�]�"���S�u��u��u����M���� S�u��u��u��M���e�[��^�É�U��WVS�u��1��ҋM�}t��$tn��C��1t]��2t1�[^_���   �%A�.�AC<.t�C���0A�f�A �   ���0��B�<	w��C��B�A<	v��f�A ����    뭍C�뙐U���E����������ES��@�]�M�uA���t�v B<$t3���u�������E��@t���t�v B<$t���u�� �1�[�Ív ���t͉�<$t�B�A��u��B븐U����u�E�u�E��E�PP�   �É�U���j �u�u�u�u�W  �ÐU���j�u�u�u�u�;  �ÐU��WVS��(�}W�u�������1҅�t
�e�[^��_�Ã��u�������1҅�u�1�;}m���E�P�U�RSV��  �E����������E����@��  �U��E�������E��@��  ��������E��@��  �E�������E��@�)  C;|�P�6�6�U�r�2�w�7�F P�5���@���   �� 9}^�ҍ�   ��   ��Q���   �f������   ���   ������   ��   ��Q���   �9������   �����      ���u�/}������   �D���$��  [����   �t��������}�f�E޴f�E��m��]��mދU؋F��9�~�V�ЋU��m��]��mދU�9�~�V�   �g�����Q�(����b�����Q�����'������   ����u-���u�|�����   ���$�P  X���   �4��1��렃�P蒸�����Ő������������먐�U��O�����U��S���]S�u�K��XZS�u�]��K���u�u�E�P�E�P�]������]���U����u�uh�u�2   ��U����u�uh�u�   ��U����u�uh�u�   ��U��WVS��  �]S�uV�������������������Ҹ�����	  P�E�phv������脟���U�B����u��6Ph�O�������a����U�B����u��6Ph�O�������>����E���@�\$�@�\$�@�\$�@�$h0v������������u�   ��������01�8��v  ���[  �U�� 1��������v ����������0����9��  �� ���P������PW�u�H  �U�ËB����t�8 u	��t[�; tV݅����݅ ����������ـ�E��@uG���$��x���hEvV�����4$�܅���ۉ�tPVhNv�������4����� G�W�����6����������������hEv��x���R赡����x����$臅��������� ���hEv�����V芡����V�a�����Y��tPV��x���RhKv������豝���x�����6�ۃ��������7����   �e�[^_�Ã��u��  ������������^_PS���������o���U��VS���]�U;�M�u~$��jQ����Y[jV������6�e�[^�Ív ���E�PPVQR�C P�$/�����   �E���ԉ�U��S���E�P�E�P�u�u����j�u��u��u���F���� j�u��u��u�F���؋]��É�U��S���E�P�E�P�u�u�>���j �u��u��u���tF���� j �u��u��u�aF���؋]��É�U��VS���E�P�E�P�u�u�]�����S�u��u��u���)F���� S�u��u��u�F���e�[��^�É�U��S���]S�u�   �E�C�]�1���U��S���]S�u�y   ǃ�       ǃ�       �    �C    �C    �C    �C    �C    �C    ǃ�   ������ �$�8*��1��]��ÐU����u�u�   1��Ív U��SP�E���]t%��P�Dw���C�$�  X�s��y��1��]��Ð��6�ԐU����u,�u(�u$�u �u�u�u�u�u�u�   1��Ív U��S���],�E�[�E�[�E�[�E$�[�u��v���C�$�  X�s�zy��1��]��Ív U����u�   1��É�U��VS�u�F����   �F��u~���~A1�9�}�����   ����uSC9�|�����   �t���X���   �h���ǆ�       ���F ��P�&���    ǆ�       �e�[1�^�É���P�+������띃�P�����F    ���j�����P�����F    ���K���U��WVS��$�}�u�w1��������;})�u���E�PVSW�X����uP�E�P�u�VC������ ;|ۍe�[^1�_�ÐU��E� �É�U��WVS���E�0���������   ���uh ��t���Y�u����1ۍ�    �$蚰����9��}	���C9�|�h��jVW�����XZ�u�5�1�������9�}/��E�P�E�P�4�h ������uP�E�P�E�PC�Q����� 9�|҃�h �����1��e�[^_�Ív U��S��<�]�SS�E�P�E�P�E�0h ��*����SS�E�P�E�P�E�0h ��*���E��E������� ��Eu���ظ�����]��Ð��������Eu	�   ���1���U��S���]�S�ԙ���$�ܗ���$蔚����� ����t�v <
tB���u��ȋ]��É�� �됐�U��E�@     �@$    �@(    �Ív U��WVS���M����   �U����   ��j�u�<����ǃ��������tA1�P�E)�P�>P�u詛��������xƅ�~w;u|ي<0t<<1t��W�~���������e�[^_���u�E�uHP�GP�1  �É<$�S�������1�N9�};]}�v �D;�U�C9�};]|��W�#������;u}����냸����딐U��WVS���M�ɋ}t]��xY��jW�^����E�U���Ҹ����tAW�u�W�u�G  ����~9�~{Vj�E�P�u�E�0�1�����Ht���u�蜮��������e�[^_�Ív 1�����S)�P�E�P�u�����������xƅ�~9�|ك��u��V���F���۸����x���뮉�Pj�E�P�u�E�1贕����Hu�1�P��)�P�E��P�u蘕��������xƅ�~�9�|�랍v U��WVS���}���ut]��xYPj�E�P�u�E�0�V�����H�����t�e�[^��_�Ð1ۉ�P��)�P�;P�u�*�������~�9�|��x	9�Stǉ������뾐U��WVS��\�E���}��   �E����   �E���#  ���  W�}���v�$f�E����vf�E����m��]��m�j�u�V菬���Ã��۸����tE���E�P�����j8h�v�Mj��M��M��EQ�E��u��]��!����� ��t��S�ͬ��������e�[^_�Ã�j�E�P薓������t5��u��S蝬���M��$覘��������Ã�S肬���E��$苘���+u�9�/1�9�}��M�
B9�|��S�Q����E��$�Z������w�����S�6����1��e����U��WVS��L�]�ۋu�}��   ����   ����   �E����   ���E�P�������j8�Eh�v�E��E�P�u��]��}��ݔ�����Ҹ����t�e�[^_�Ã�j�E�P�����]+]�����v���t���E�P�J����������;]u���E�P�2�����믉�1�멸����뢐U��U���t<
tB���u��Ív � ��U��U��J��S�M�]~����ACJ���[��U���j4�u�u������Ð��U��SP�]�ۋE�p���� t��t��Ph���������؋]���U��p��É�U�����É�U���p�    ��� �Ð�U��WVS��   �}�E�  W��  ����u�����e�[^_�Ð��W�  �����P  ��W�  ����u1��σ�W�  �����  ����d���VW�(  ����uD�E�8 ��  ��d�����  ��HP��d���hw��h���S�o���YXS�u��������VW�G  ����uD�E�8 �`  ��d����I  ��HP��d���hw��h���S����XZS�u诓������VW�f  ����uD�E�8 ��  ��d�����  ��HP��d���h%w��h���S�Ŕ��YXS�u�Z�������VW�e  ����uD�E�8 �v  ��d����_  ��HP��d���h.w��h���S�p���XZS�u��������VW�d  ����uD�E�8 �  ��d�����   ��HP��d���h8w��h���S����ZYS�u谒��������X���PW�]  ���������E�8 ��   ��VW�  ����t
ǅd���    ݅X�������������E����@uG��d�����u=��6P��\�����X�����d���hDw��h���S������S�u������������H����hdP��������h�����6������hdP�֑�����������6������hdP趑�����t�����6�'�����hdP薑�����������6������hdP�v�����������6�=�����hdP�V�����������hRw�u�>����������������d���VW��  ������  ��VW�_  ����u'�E�8 ��  ����d����4�|��u����������d���PW�  ����uB�E�8 �4  Q��d���h�s��h���S����XZS�u蛐���<$��  ������  ����d���PW�  ����u2�E�8 ��  P��d���haw��h���S譑��^XS�u�B���������d���PW�  ����u2�E�8 �N  Q��d���haw��h���S�d���XZS�u�����������X���PW�  ����ub�E�8 ��   ����d���PW��  ����t
ǅd���    ����\�����X�����d���hTw��h���S������S�u耏��������d���PW�  ����������E�8 ucP��T���P��P���P��d����  X��d�����T�������P���x+��YPh[w��h���S�r�����S�u�������z����Rw�Ӄ�hdP������늃�h
;P�֎�����������h
;P�������������hdP誎�����=�����hfw�u蒎����������hdP�|�����������hdP�f������b���Q��d���h�s��h���S規��XZS�u�;������������U��VS���]�uS��  ����t9��SV�C  ����t�e�[1�^�Ív �E�w�E�����e�[^������v ��SV�   ����u��E�w�E�����эv U��WVS��X  �������ES�}ǅ����    ǅ����    ǅ����    ǅ����    �������l  ��1҅�u�e�[^��_�ÐP������P������PS�#  ������  ��������VS�  ��1҅�t���������PV��  ��1҅�t�P������P������PS��  ��1҅�t���S�  �����   tǅ����   ���S�  ��1҅��O�����������VjjW�  �� 1҅��.����   9�   ǅ����   <���w)�$�<x��������W�e  ��1҅������������B9�������~ŋ�������u2��������u
�   ������������W�  ��1҅�������؃�W�T  ������������W�`  녃�������W��  �q�����������W�  �]�����������W�C  �I���Q������������W�  �1�������S�  ����������t�������   ������������������PS�  ����tӋ�������������������P������P�  ��1҅��   �����P������P������PS��  ��1҅��������S�"  ����t
ǅ����   P������P������PS�  ����������������8:�   �����@V������������P������PS�i  ��1҅�����������t1��	����������8:�   tM��������PS�  �����y�����������P������P��  ��1҅������ǅ����   �G���@������������P������P������PS�A  ��1҅��}����������`����   �m����U��WVS��X�]�S��E�]��E�    �E�    �E�    �E�    �E�    �E�    �E��  �Ẻ$�v  1���1҅��   ��   �����E�P�E�P�E�P�E�PS�  �� ����   �E�9�~��9�}�ǃ�t�U����   ��w��$�Xx�}�f�Eִf�E��E��m��]��m���}�f�Eִf�E��E��m��]��m��x����}�f�Eִf�E��E��m��]��m��Z����}�f�Eִf�E��E��m��]��m��<����}�f�Eִf�E��E��m��]��m������E؋E��]��E�����1ҍe�[^��_�Ã�S�X  ��1҅�u���u�WVj�u�  �� 1҅�u�9����u��0��w!�$�tx���u��u�  ��1҅�u��E�@9��E��~ЋE̅�u�   뀃��u�<  ������u��u�I  뼃��u��u�  묃��u��u��  뜃��u��u�5  �P�u��u��u�  �x����v U��U1��� t��	t
��
t�Ív �   ���U��E��0<	�����ÐU��VS�u����P��������t�C���e�[^�ÐU��WVS���u�    �u�}�����E����    ����P��������t��������DЉC��֋��~�U������e�[^��_�Ív U��WVS��  �u�L����E�0�E�     �������E���     �����P�
�������t��EFG� ����.t6Q� �uh�O������P������1�Ht
�e�[^��_�ËE�0�   ���.FG�����P��������t���EFG� ��U��VS�]����   tA����V�U��������   u)�E��t.���C�P�Y����É4$�O���1҃�9���e�[��^�Ív 1���U��WVS���u�}�4����E�0���E�    ����t,����S���������u��S�&   �FG���E�   ��� �E�0�E��e�[^_�Ív U��U�B�<w�� ���Ív U��WVS���}1۾������4�W�p�������tC��~�1��e�[^_�ËE�S��   ���U��S��  �]�������������P������P������1҅�t������bu������cu	������ t	1҉Ћ]��Ë�������   ��U��WVS���]�E�    �<+t<-�E�   t1ҍe�[^��_�Ã��sV�������1҅�t����{W������1҅�tʃ��CP�E�������1҅�t����[S������1҅�t�����������M�F���P�M���0����ɋU�t�؉�   �\�����U��WVS��  �U��u�u�u������S���������������u1��e�[^_�Ív ��������PS��������t܍�������y�   ��t�������x�   �u�U�   �������U��   뚍������!z�   ��t:�������x�   �t&��������mu&������ou������nu������ u�E�    딀�du������au������yu	������ t�������x�   ��u�U�   �Q����������wz�   ��t�������#x�   �u�E�    ������������z�   ��t4�������)x�   �t ��mu)������iu ������nu������ u�U�   �������������z�   ��tD�������1x�   �t0��s�;���������e�.���������c�!��������� �����E�    �\����v U��S���]S��������8-t
1��]��Ív @��   ���U��S�� �]�S�E�E������E��$PP�E�PS�x����� �������]���U��S���]S��������8 �����]��ÐU��E�@,�������ÐU��E�P,�������ÐU��E�@,   �ÐU��E�@,    �ÐU��U1��z, ���B,��U��S���]�E��E�C�E�C�E�C�C    �C    �C    �C    �C     �C$    �C(    S��  �C,   ���]�]���J   ��U��M��E��Q�E��Q�E��Q�E���   �U����u�   ���������ÐU��SS�]�H��v��h�xj��y����]���Qjj�s�	  ����u��h�xj���Rjj�s��  ������   �S;S��   ���t6Ht�{t1�룋C��y���h�xj�닐�{t܃�h yj��u�����R�r   ����t���s�`   ����t(���s�b   ����u�뒃��s�L   ����u��h`yj���������h�xj�������h�xj��������U���jj�u�  ��U���jj�u��  ��U��E�8�����Ív U��E�8�����Ð��U����E�p�p�u�  �Ív U��VS���]�uS��������tU��Sj��������t3��V�   ����t	�e�[1�^���E�y�E�����e�[^�������E�y�E�������E�y�E������U��S���]�s0S�m���������u�S0�E��ȋ]��ÐU��VS���]S�uV�?�������u�^0�e�[^�É�U��E�@0�����1�Ív U��E�  =�  ������U��WVS��d�E�P�}W�]�g�������t�e�[^_�Ã�S��������u��h�yj�������׍v ��j jjj�u�V�\����� +]�x��SV�b  XZVW��  룃�V�"���YX����U���j �u�d����É�U��M��Sx�Ȼ<   ����ыU��E��$�É�����U����E�p�p�u��  �Ív U��VS���]�uSj���������t?��x��S��������t��~�e�[1�^�É��E�y�E�����e�[^�������v �E�y�E������U��VS���]�uSj�b�������t_��x?��S�>�������t�F���w'��S�:�������t�{t���e�[1�^�Ív �Ez�E�����e�[^��?����v �E'z�E������U��VS���]Sj�u���������t��xg��S��������u1��e�[^�É����E�PS�c  ����u���E�PS��  ����uσ�S��������~RP�u��u��  ��9�~���h=zj�����뚍v ��hRzj���U��VS���]�uSj�.�������t7��x�{t���e�[1�^�Ív �Efz�E�����e�[^��3����v �E|z�E������U��VS���]�uSj���������t7��x�{t��;�e�[1�^�Ív �E�z�E�����e�[^�������v �E�y�E������U��S���E�]�]�Sj�d�������tI���E���������Et!�{t��m�E�������t	1��]��É��E�z�E�����]���U�����E�z�E������U��S���]�uj���������t%��x1��]����E�z�E�����]�������v �E�z�E������U��S���]�sS����������u�S�E��ȋ]��ÐU��WVS���}W�uV����������t�e��[^_�Ív ���~V�@�������t��F    ��U��S���]�sS����������u�S�E��ȋ]��ÐU��WVS���}W�uV����������t�e��[^_�Ív ���~V���������t��F    ��U��S���]�sS�����������u�S�E��ȋ]��ÐU��VS���]S�uV��������u�^�e�[^�É�U��S���]�sS�!���������u�S�E��ȋ]��ÐU��VS���]S�uV���������u�^�e�[^�É�U��S���]�s S�1���������u�S �E��ȋ]��ÐU��VS���]S�uV��������u�^ �e�[^�É�U��VSQ�u�v(�v$V�?���������u�V$�N(�E��H�e���[^�Ív U��WVS���uV�]S�}W��������u�_$�w(�e�[^_�ÐU��S���]�sS�Q���������u�S�E��ȋ]��ÐU��VS���]S�uV�#�������u�^�e�[^�Ð�U��M�U9�S�E1�9�	9��   �؋$�Ð1�9��9��琐U��SR�]�;��t�C,��u���]��Ív �؃��s�{�������t��v�{�C���{� {�{���{���({�{ ���0{�{$���U��WVS��T�uV�u��
  �����h  �E�8�  �}�O,���  �F,����   �����   ����   ����   ��u[�^��?PjVW�1
  ���E�8t
1��e�[^_��j��p�pW�b  Y[W�u��������؉�PSVWK��   �����뭋^��PjVW��   �PSVWK��	  ��������^;^|�PSVWK�   ��;^}��s�������@������@����^;^�V���PSVWK�z	  ��;^}��?�����F,������P�]�S�G���Z�U�r�����������j��U���r�D PS�  �߃������v �[����������U��WVS��\  �u����}�]��  Ht�e�[^1�_�Ív ��W��(���Pǅ����    ��������w��$�@{�F$�G$������EuT������ٽ������f�������5�m�f��������٭����۝����٭�����������R����P�$�V$���G$����������^$�T���Q������j��H�����(���PV�������0����F�W9�~
)ЉF������������PV�
  Y�F,������������x���������   �^�FKH�ۉ� ���~P�v,S�v�
  K� ��������F������F ������F$�V(������G+F��@�FV����������F   �F   �F     �F    �F$    �F(    Y[������SV���������FH�������G+F@���FV������F   XZǅ����    ������R뼋^�G9�)��)ٸ���*�������)�@�������@���F�ËG������)Å��^�����S������j��(�����8���S�r����V�G9�~')��������V�����������P��<���j�:�����V������R�P���j�jj������S�	  ��������PS�B  �^��;_ǅ����   ~
�^�ڋG�Pj������P������R���������������������������  ���������;_~�봋^�G9�}+)؍H�����*�������)�@�������@�ÉF�ËG)Ë��������^�����P������j��@����K����N �G 9�}%)�H�<   �ә��@�������@�����F ���G ������)��҉N �N�����������D���Pj��(���R�������V��h���Pǅ����    �����XZW�U�R��������������$�\{�F$�G$������E������   ��ٽ����f���������f������٭����ە����٭����������P�$������E����@ug�����������5�m��٭����۝����٭�����������R����P�$�V$���G$����������^$�K���Q������j�]ȍE���������������5�m�8{٭����۝����٭���������뫋V�G9�|
)V�����)Ѓ��FV�|���ǅx���    �F    _X��h��������^�G9�}*)؍H�����*�������)�@�������@���F�ËG)Ë��������^�����������P�]�j�2����V�G9�|
)V�]���)Ѓ��FV������E�    �F    �F     �F$    �F(    �Q����^�G9�}+)؍H�����*�������)�@�������@�ÉF�ËG)Ë��������^�����P������j�]������N �G 9�}%)�H�<   �ә��@�������@�����F ���G ������)��҉N ������������E�Pj�U��?����U��WVS���]�C�S9ЉE����U�~:��~5��m�v ���  ����  ���o  I;M��^  ����؋E���E  �C,���:  �3���%  �}���   Nt4�M��u�;t
�e�[^1�_�ËC��x	�C,   ���؉C�C,    �؃}�~�V�s,�s�s�  ��9C~�W�s,�s�s�z  )C�C����t@�C�ƋC@���Cu�C   �C   뫃}��d�����t1�K���S�������*��׉�����)Ǎ��)�{�K�.����C���E�������I����*�������)ϋC����Cu�C   ���)E�U�S������[��������3������������s�����������*��׉�����)Ǎ��)�{�s�_������V����C$������u8�}�f�E����f�E����m��]��m�}�����{ P�$$���[$�����������s ��;�������<   ���C�@����)Ɖs �����U����E���U�Mw�$�x{�A$�B$�Z$�:t��j R�d�����1��Ð��j��AB�ًAB�ыAB�ɋAB���A B 빐U����u�u�   ���������É�U��VS���]�uS���������   u�e�[��^�Ív ��V���������   t߃�V�����������   �C9Fs��P��������t���v��������tA���s��������u1�닃��v�x�������u��E�{�E�����e�[^������E�{�E�������E�{�E�������E |�E������U��WVS���E�U�]�u�E��}�U�S��������tQ�   �C����C�U�S���������u�C�U���e�[^1�_�Ã��s�������������D �Սe�[^_��<���U��E���$P�E�P�E�P�E�P�u�Z����� ��t�����Ã��u��u��u��u��u�q����吐�U��VSS�M�ɋUtD1���t71���x11���   u�d   �ȉ֙����u��  �ȉ֙����u�   ��Z[^�É��E@|�E����Y[^��Q����U����E���Uu�E�|�E������,�����RP�f�����������m  ��U��SP�]�C����M�Uw.��t�����Ћ]��Ív ��RQ���������   u����E�|�E�����]�������U��WVS��   �uV�}��������������u�e�[^��_�É���j W�u�6�E�P� ����� �������uԋF��`�����`����E9ÉF}*��m����#  ����  ����  C;]|��؋V9���   �E����   ��V�����������V��1�9���T�����~'����w�$��|��T���9Ft�   K��u9�ۅ�tXVWW��h���P�  XZ��h���PVǅx���   ǅ|���   �E�   �E�   �E�   �E�    �E�  �?�������]����   �V�];�`���}����w�$�}�F    �C;�`���|�9׉�~���w�$�(}�F    �K9����F    �~1��e����F    ���F    ���F    ���F     ���F$    �F(    ��F    ��F    �x����F    �l����F     �`����F$    �F(    �M�����V�(���������   ǅd���    �V9���������d������d�������\���VSS��h���P�0  �F��x����F��|�����\���F�E��F�V(�E��F �E��F$�U�ZY�E���h���PV�;�����d�������~	���}���K9���s������v,�v�m�������d����L�����T���9F������F��������F �������F$����������E��@�����������F�@��F�F    �/�����t ���!������N �F$�^$�F     �
����F�@����F �F    ������F�@��F�F    �����U��VS���]�uj �u�ujV������S��������u
�e�[^�Ív ��S�'�������t�u�e�[^��6�����U��VS�6`���H�-H���1�9�s�Ɛ��H�C9�r�[^��U��SP�H�-H������X�u�]���6   ����H���K��u���U��SR�������t���Ћ���u�X[��U��SR�    [�ê_  �e���]���                                                          GRASS GNU GPL licensed Software Sample semivariogram of a GRASS sites list.                     basename of a graphing data/commands files (implies -p)         which decimal attribute (if multiple)                           lag tolerance must be less than half nominal lag                error scanning anglular tolerance                               No sites found. Check your region.                              I'm really not smart enough to deal with your projection        Computing sample semivariogram ...                              Plotting ...                                                    Ran out of memory; try reducing your region size                Decimal attribute field 0 doesn't exist. sites name of a sites file old,site_lists,sites,input nominal lag distance lagtol direction direction of semivariogram angtol direction tolerance graph 1 Quiet Plot sample semivariogram GRASS_GNUPLOT error scanning lag error scanning lag tolerance error scanning angle  site_lists %d sites found
 %g %g %d
 Some pairs of data ignored oops, not enough bins can't open sites file [%s] sites file [%s] not found             �?�cܥL@                                        out of memory
                                                  plot %s.gp %s.dat Error opening temporary file                                                       �v@                        set title 'Sample Semivariogram'
                               plot %s using 1:2 title "" with %s
                             plot '%s' using 1:2 title %c%c with points%s                    Saving plot files ...                                           Unable to open the temporary file. #h g N(n) 
 cd ' set size 1,0.9
 set nokey
 set xlabel 'lag (h)'
 dots points %s %s                                          G_malloc: out of memory G_calloc: out of memory G_realloc: out of memory                        G_distance_point_to_line_segment: shouldn't happen
              code=%d P=(%f,%f) S=(%f,%f)(%f,%f)
          �                -------------------------------------
 ERROR libgis %s:  WARNING %s: GRASS_STDERR %s/GIS_ERROR_LOG program: %-10s %s
 user: cwd: date: error: warning: mail '%s' GIS %s: %s
 
%*s                                                                                     �?-DT�!	@     �f@      @       �      �?                invalid a: field %s in file %s in %s                            invalid ellipsoid %s in file %s in %s                           invalid es: field %s in file %s in %s                           No ellipsoid info given in file %s in %s                        Line%s%s of ellipsoid table file <%s> %s invalid                unable to open ellipsoid table file: %s PERMANENT PROJ_INFO ellps sphere proj Unable to open file %s in %s a=%lf e=%lf f=1/%lf b=%lf %s/etc/ellipse.table %s  "%32[^"]" %s %s  %d are           region for current mapset %s
run "g.region" DEFAULT_WIND default region %s is invalid
%s                                                                        GISBASE                         ERROR: System not initialized. Programmer forgot to call G_gisinit()
 @(#) 5.0.3 (October 2003) MAPSET %s not found MAPSET %s - permission denied              unable to determine user's home directory cd; pwd                                                                                                               Illegal filename.  Cannot be '.' or 'NULL'
                     Illegal filename. character <%c> not allowed.        /locale    LOCATION  << %s >>  not available LOCATION_NAME %s/%s                                           MAPSET is not set MAPSET        can't make mapset element %s (%s) mkdir                                                         SEARCH_PATH                                                     %s %s %s %s@%s                  EmbedGivenNulls: wrong data type!                               Null values have not been initialized.                          G_gisinit() must be called first.                               Please advise GRASS developers of this error.
                  G_set_null_value: wrong data type!                              G_is_null_value: wrong data type!                               G__check_null_bit: can't access index %d. Size of flags is %d (bit # is %d                      G__open(w): xmapset (%s) != G_mapset() (%s)
                    G__open(r): mapset (%s) doesn't match xmapset (%s)
 r+          unable to open raster map [%s in %s]                            [%s] in mapset [%s] - in different projection than current region:
 found map [%s] in: <%s>, should be <%s>                     [%s] in mapset [%s] - in different zone [%d] than current region [%d]                           [%s] in [%s] - bytes per cell (%d) too large                    [%s] in mapset [%s]-format field in header file invalid         unable to open [%s] in [%s] since it is a reclass of [%s] in [%s] which does not exist          G__open_raster_new: too many open files                         opencell opening temp null file: no temp files available        Can't write embedded null values for map open for random access G__open_raster_new: no temp files available                     opencell: %s - illegal file name                                G_set_fp_type() can only be called with FCELL_TYPE or DCELL_TYPE                                the map %s is not xdr: byte_order: %s                           invalid type: field %s in file %s                               G_set_quant_rules can be called only for raster maps opened for reading Too many open raster files GRASS_FP_DOUBLE opencell: %s - bad mapset opencell: too many open files unable to find [%s] in [%s] fcell g3dcell cell_misc/%s f_format unable to find [%s] Unable to open %s double float byte_order %s - ** illegal name **                                Sorry <%s> is not a valid option
                               <?xml version="1.0" encoding="UTF-8"?>
                         <!DOCTYPE task SYSTEM "grass-interface.dtd">
                   	<parameter name="%s" type="%s" required="%s" multiple="%s">
   Sorry, <%c> is not a valid flag
                                Sorry, <%s> is not a valid parameter
                           
Error: Missing value for parameter <%s>
                       
Error: value <%s> out of range for parameter <%s>
             
Error: illegal range syntax for parameter <%s>
                
ERROR: Required parameter <%s> not set:
 (%s).
                
Error: option <%s> must be provided in multiples of %d
               You provided %d items:
  Programmer error: no flags or options
                          
FLAG: Set the following flag?
 
PROGRAMMER ERROR: first item in gisprompt is <%s>
                     Must be either new, old, mapset, or any
 --help --interface-description 
Usage:
  = 
Parameters:
   %*s   %s
   %*s   default: %s
 
Flags:
   -%c   %s
 [, ,...] [ 
Description:
 ?? &amp; &gt; &lt; <task name="%s">
 integer no 	</parameter>
 	<flag name="%c">
 	</flag>
 </task>
 		<description>
			 
		</description>
 		<values>
 			<value> </value>
 		</values>
 			<default>
			 
			</default>
 age element prompt 		<gisprompt  />
 %s="%s"  		<keydesc>
 			<item order="%d"> </item>
 		</keydesc>
 yes 	<description>
		 
	</description>
   %*s   options:  %s, 
 %*s 
   Sorry, <%s=> is ambiguous
        Legal range: %s
        Presented as: %s
 %d-%d %lf-%lf     %s? 
OPTION:   %s
      key: %s
 YES required: %s
 %s=%s 
You have chosen:
  %s
 Is this correct?  Sorry, %s is not accepted.
    Try again?  enter option >   options: %s
 multiple: %s
 NO   format: %s
 to accept the default +,-./:=_                                                     %4d%%                                                      -c /bin/sh                                                                                                                                                      degrees degree feet foot units unit meters meter State Plane x,y UTM Other Projection Latitude-Longitude                                                        PROJ_UNITS Unknown projection inch datum                                                                                        G_truncate_fp_map: can't write quant rules for map %s           G_quantize_fp_map: raster map %s is empty                       G_quantize_fp_map: can't read fp range for map %s               G_quantize_fp_map_range: can't write quant rules for map %s     Cannot write quant rules: map %s is integer                     Cannot write quant rules for map %s                             can't read f_range file for [%s in %s]                          G_read_range(): can't read quant rules for fp map %s@%s         can't read range file for [%s in %s]                            G_write_range(): the map is floating point!                     can't write range file for [%s in %s] f_range Too many open files %d%d%d%d %ld %ld
                                             duplicate e-w resolution field  duplicate n-s resolution field duplicate projection field duplicate zone field zone field missing nort duplicate north field sout duplicate south field east duplicate east field west duplicate west field e-w  n-s  rows duplicate rows field cols duplicate cols field form duplicate format field comp duplicate compressed field rows field missing cols field missing east field missing west field missing south field missing north field missing projection field missing %[^:]:%[^
] %d%1s line %d: <%s>              I'm finding records that do not have a floating point attributes (fields prefixed with '%').    decimal field %i not present in sites file                      Reading sites list ...                   cannot allocate memory failed to guess format          %s/%s/cell_misc/%s/reclassed_to Illegal reclass format in header file for [%s in %s]            Too many reclass categories for [%s in %s]                      Unable to create header file for [%s in %s] null reclas %[^:]:%s maps cellhd reclass
 name: %s
 mapset: %s
 0
 a+ %s@%s
 #%ld
 Illegal reclass request Illegal reclass type #%d                                                 rm -rf '%s'                     G_set_window(): projection/zone differs from that of currently open raster files G_set_window(): %s                             G_site_new_struct: invalid # dims or fields
                    
PROGRAMMER ERROR: G_site_describe() must be called
                    immediately after G_fopen_sites_old()
                  Memory error in writing timestamp                               
PROGRAMMER ERROR: G_site_get_head() must be called
            Memory error in allocating timestamp                            WARNING: %s needs modified for the new Sites API
 %[^|]|%[^|]|%*[^
] ERROR: ebuf %s nbuf %s
 %lf| #%lf #%f %s|%s| %%%s  @"%s"  @%s  #%g  #%d  #%s  . time|%s
 Illegal TimeStamp string labels|%s
 form|%s
 desc|%s
 name|%s
 name| desc| form| labels| time| %.8f site list point|%[^|]|%[^|]|%[^
] %s|%s|%s
 # %s%s%g  % @ %s%s"%s" %s%s%d       �                                                                            WARNING: can not create a new process
                                                          %d.%d /                         Invalid timestamp specified for %s map %s in mapset %s          Can't create timestamp file for %s map %s in mapset %s          Invalid timestamp file for %s map %s in mapset %s               Can't open timestamp file for %s map %s in mapset %s %s / %s cell_misc timestamp raster dig_misc vector grid3                                                                                                                                                                                                                        �V@     �V�     �f�%lf%1s                                                                                                                                  (y/n)  [n]  [y]                                                 North must be larger than South North must be north of South Invalid coordinates East must be larger than West Illegal latitude for South Illegal latitude for North Illegal e-w resolution value Illegal col value Illegal n-s resolution value Illegal row value                                                                                              Enter 'list' for a list of existing %s files
                   
** %s exists. ok to overwrite?                                 
** %s - exists, select another name **
                        Enter the name of an existing %s file to cancel request Enter %s file name 
%s
 Enter 'list -f' for  an extended list Hit RETURN %s
 <%s>
 ** illegal request **
 
** %s - not found **
 
** %s - illegal request **
 
**<%s> illegal name **
 a list %s Enter a new %s file name ask: can't happen %s%s%s%s    ��x�M�U�a�                            Unable to open automatic MASK file MASK                                                         closecell: can't move %s
to cell file %s                        Error writing floating point format file for map %s             closecell: can't move %s
to null file %s                        Can't write f_format file for CELL maps  can't write quant file! f_quant mv %s %s xdr lzw_compression_bits                                                                                      GISRC GISRC - variable not set %s not set                                                                                                                                                       Fail of initial read of compressed file [%s in %s]              Can't read header file for [%s in %s]
                          It is a reclass of [%s in %s] whose header file is invalid
     It is a reclass of [%s in %s]   whose header file can't be opened                               Can't open header file for [%s in %s] Invalid format
 which is missing                                                                                          GISDBASE                        Histogram for [%s in %s] missing (run r.support)                Invalid histogram file for [%s in %s]                           Can't read histogram for [%s in %s]                             can't create histogram for [%s in %s] histogram %ld:%ld %ld:%ld
                                can't get history information for [%s] in mapset [%s]           can't write history information for [%s] hist generated by %s                                   G_random_d_initialize_0: write failed in row %d.
               G_random_d_initialize_0: xdr_double failed for index %d.
       G_random_f_initialize_0: write failed in row %d.
               G_random_f_initialize_0: xdr_float failed for index %d.
                                                                                                        ----------------------------------------------
                 %s files available in mapset %s:
 hit RETURN to continue --> no %s files available
 $GRASS_PAGER ls %s 
%-18s %-.60s
 ls -C %s                                  dd:mm:ss{N|S} ddd:mm:ss{E|W} dd:mm:ss 0%f %d:%02d:%s%c %d:%02d%c %d%c 0       N@      $@                                        sn we %se %d:%d:%d.%[0123456789]%[^
] %d:%d:%d%[^
]     �������?      �@                                                        Unable to create header file for [%s]                           %s: %s is not integer! Use G_put_[f/d_]raster_row()!            %s: map [%s] not open for random write - request ignored        %s: unopened file descriptor - request ignored                  %s: map [%s] not open for write - request ignored               %s: map [%s] not open for sequential write - request ignored    map [%s] - unable to write row %d                               xdr_double failed for index %d of row %d.
                      xdr_float failed for index %d of row %d.
                       unable to find a temporary null file %s                         G__open_null_new(): too many open files!                        can't put float row into integer map                            can't put double row into integer map G_put_map_row G_put_map_row_random G__put_null_value_row G_put_raster_row error writing null row %d
                      The floating data range for %s@%s is empty                      The integer data range for %s@%s is empty                       G__quant_import: attempt to open quantization table for CELL_TYPE file [%s] in mapset {%s]      quantization file in quant2 for [%s] in mapset [%s] is empty    quantization file [%s] in mapset [%s] %s quant2/%s empty truncate round %lf:%lf:%d:%d *:%lf:%d %lf:*:%d *:%.20g:%d
 %.20g:*:%d
 %.20g:%.20g:%d                                                  colr colr2/%s                                                   proj:       %d
 zone:       %d
 north:      %s
 south:      %s
 east:       %s
 west:       %s
 cols:       %d
 rows:       %d
 e-w resol:  %s
 n-s resol:  %s
 format:     %d
 compressed: %d
                                                                                                 category support for [%s] in mapset [%s] %s                     category support for vector file [%s] in mapset [%s] %s invalid dig_cats dig # %ld %lf:%lf:%[^
] %d:%[^
] %f %f %f %f no data # %ld categories
 %.2f %.2f %.2f %.2f
 %.10f %s:%s:%s
                                                                            1.1.4   )\���(�?      (@                                        Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec %d year%s %d month%s %d day%s %d hour%s %d minute%s %.*f second%s - %02.*f %s%02d%02d  bc                       Invalid interval datetime format                                Invalid absolute datetime format jan feb mar apr may jun jul aug sep oct nov dec years months days hours minutes seconds    n	L	�	�	�	�	
X����:�����invalid datetime 'mode' invalid datetime 'from' invalid datetime 'fracsec' invalid datetime 'from-to' invalid datetime 'to'                     invalid absolute datetime 'from'                                invalid relative datetime 'from-to' invalid datetime timezone datetime has no minute datetime not absolute                           invalid datetime year datetime has no year invalid datetime month datetime has no month invalid datetime day datetime has no day invalid datetime hour datetime has no hour invalid datetime minute invalid datetime second datetime has no second invalid datetime fracsec datetime has no fracsec                     �v@     �@     A    ~~A      �?�!_"~#�#�$�$�!�!�&�&'h'�'�%�*�*�*�*�*�*�*            illegal datetime increment interval                             datetime increment too precise  datetime increment mode not relative                            datetime_is_leap_year(): illegal year                           datetime_days_in_year(): illegal year                           datetime_days_in_month(): illegal month         �.�.�.�0�0�0�0T/L/�/�/�/�/�/x/p/�/�/�/�/�/                                    ��2�2�2�2�2�2    �2          �?�2               �2�2�2    ����H=�2   �2�2�2�>    �2    �2�2�2�2�2   �2�2        �2�2    �2�2              �2                    -x �2�����2�2�O�2�2                    �2                            �Q      �?�Q      �?�Q����ׁ�?^R�
F%u�?            �2�2�2�2�2�2�2�Y�2�2�2    �2�2�2�2    �2�2�2    �2�2�2�2�2�2�2�2         �2            �2�2@   �2�2�2                        �2�2�2�2�2    �2�2�2�2�2�2�2�2    �2�2�2�2                        �2                           t��� �\�t������t��2�2�2�2�2�2�2�6�2�2�2                �v�v�v�v�v�v�v�v wwww                �w�w�w�w�w�w�w�wxx	xx                                                             ;      �       �   h2   (�   ��   P�
   J                  �   �           X�   8�             ���o؎���o   ���o
�                                                ����    ����        0�        N�^�n�~���������Βޒ�����.�>�N�^�n�~���������Γޓ�����.�>�N�^�n�~���������Δޔ�����.�>�N�^�n�~���������Εޕ�����.�>�N�^�n�~���������Ζޖ�����.�>�N�^�n�~���������Η                     GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  GCC: (GNU) 3.2.2 20030222 (Red Hat Linux 3.2.2-5)  .shstrtab .interp .note.ABI-tag .hash .dynsym .dynstr .gnu.version .gnu.version_r .rel.dyn .rel.plt .init .text .fini .rodata .eh_frame .data .dynamic .ctors .dtors .jcr .got .bss .comment                                                     ��                              �                     !         (�(  (               '         P�P  p              /         ���
  J                 7   ���o   
�
  �                D   ���o   ؎�  `                S   	      8�8                   \   	      X�X  �              e          �                     `         8�8  �                k         ؗ�  ��                q         h2h�                   w         �2�� �J                           D}D�                   �         `�`� �                  �         0�0 �                �         �                   �         �                   �         �                   �         � t                �         ��� L\                 �              � O                               � �                  